ClockSynthesizer.vhd