-- $Id
-- This package contains constants used by the cic_v1_0

package cic_pack_v3_0 is
  constant c_interpolating_filter: integer := 1;
  constant c_decimating_filter   : integer := 2;
  
  constant programmable : integer := 1;
  constant fixed        : integer := 2;
end cic_pack_v3_0;
  
