-------------------------------------------------------------------------------
-- DESCRIPTION: 
--
-- NOTES:
--
-- $Author$
-- $Date$
-- $Name$
-- $Revision$
--
-------------------------------------------------------------------------------

---------------
-- LIBRARIES --
---------------

library ieee;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

----------------------------------
-- COMPONENT PACKAGE DEFINITION --
----------------------------------

package uSoCControllerPackage is

  -- CONSTANTS

  -- TYPES

end uSoCControllerPackage;

-------------------------------------------------------------------------------
-- $Log$
-------------------------------------------------------------------------------
   
