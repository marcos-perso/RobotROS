-------------------------------------------------------------------------------
-- DESCRIPTION: 
--
-- NOTES:
--
-- $Author$
-- $Date$
-- $Name$
-- $Revision$
--
-------------------------------------------------------------------------------

---------------
-- LIBRARIES --
---------------

library ieee;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

----------------------------------
-- COMPONENT PACKAGE DEFINITION --
----------------------------------

package PWMGeneratorPackage is

  -- CONSTANTS
  constant C_PWMCOUNTER_MAX : integer := 64000;
  constant C_NB_BITS_PWM_COUNTER : integer := 24;

  -- TYPES

end PWMGeneratorPackage;

-------------------------------------------------------------------------------
-- $Log$
-------------------------------------------------------------------------------
   
