DualRAM_8x32.vhd