RAM1024x32.vhd