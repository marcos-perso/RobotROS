--------------------------------------------------------------------------------
--This file contains code that has been derived from code licensed to
--Xilinx by QinetiQ ltd.
--------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /   Vendor: Xilinx
-- \   \   \/    Version: 1.0
--  \   \        Filename: $RCSfile: floating_point_v1_0_xst.vhd,v $           
--  /   /        Date Last Modified: $Date: 2010-07-10 21:43:11 $ 
-- /___/   /\    Date Created: Dec 2005
-- \   \  /  \
--  \___\/\___\
-- 
--Device  : All
--Library : xilinxcorelib.floating_point_v1_0
--Purpose : Floating-point operator behavioral model
--Revision History:
--   16 Feb 05 : Added assert statement to catch unsupported C_OPTIMIZATION.
--   28 Feb 05 : Removed non static array definition i.e. (ew=>'1', others=>'0')
--               from fpMul, fpDiv and fpSqrt. Changed all architectures to
--               behavioral.
--    1 Mar 05 : Added functions to support multiplier type.
--   14 Mar 05 : Detected sign of zeros in fpAdd to get -0+-0 =-0.
--               Correctly signed zero when underflow.
--   16 Mar 05 : Removed underflow in fpMul when one input is zero. It now never
--               signals an underflow when one or both of the inputs are zero.
--               Added divide by zero exception to divider when a finite,
--               non-zero number is divided by zero. 
--   22 Mar 05 : Infinity divided by zero does not raise a divide by zero
--               exception.
--   28 Mar 05 : Modified RDY output to get correct behavior with STATUS_EARLY.
--   21 Apr 05 : Included SCLR on new_operation in order to reset RDY signal
--               correctly. Use undelayed operation for start detection.
--               Added SCLR to input delays so that output is set to zero 
--               (i.e. 0+0=0).
--
--------------------------------------------------------------------------------    
--  Copyright(C) 2005 by Xilinx, Inc. All rights reserved.
--  This text/file contains proprietary, confidential
--  information of Xilinx, Inc., is distributed under license
--  from Xilinx, Inc., and may be used, copied and/or
--  disclosed only pursuant to the terms of a valid license
--  agreement with Xilinx, Inc.  Xilinx hereby grants you
--  a license to use this text/file solely for design, simulation,
--  implementation and creation of design files limited
--  to Xilinx devices or technologies. Use with non-Xilinx
--  devices or technologies is expressly prohibited and
--  immediately terminates your license unless covered by
--  a separate agreement.
--
--  Xilinx is providing this design, code, or information
--  "as is" solely for use in developing programs and
--  solutions for Xilinx devices.  By providing this design,
--  code, or information as one possible implementation of
--  this feature, application or standard, Xilinx is making no
--  representation that this implementation is free from any
--  claims of infringement.  You are responsible for
--  obtaining any rights you may require for your implementation.
--  Xilinx expressly disclaims any warranty whatsoever with
--  respect to the adequacy of the implementation, including
--  but not limited to any warranties or representations that this
--  implementation is free from claims of infringement, implied
--  warranties of merchantability or fitness for a particular
--  purpose.
--
--  Xilinx products are not intended for use in life support
--  appliances, devices, or systems. Use in such applications are
--  expressly prohibited.
--
--  This copyright and support notice must be retained as part
--  of this text at all times. (c) Copyright 1995-2005 Xilinx, Inc.
--  All rights reserved.
--
--------------------------------------------------------------------------------

LIBRARY IEEE;USE IEEE.STD_LOGIC_1164.ALL;USE IEEE.STD_LOGIC_ARITH.ALL;LIBRARY XILINXCORELIB;USE XILINXCORELIB.
FLOATING_POINT_V1_0_CONSTS.ALL;USE XILINXCORELIB.FLOATING_POINT_PKG_V1_0.ALL;ENTITY FLT_PT_OPERATOR IS GENERIC(C_FAMILY:STRING;
C_WIDTH:INTEGER;C_FRACTION_WIDTH:INTEGER;C_OPTIMIZATION:INTEGER;C_MULT_USAGE:INTEGER;C_HAS_STATUS:INTEGER;C_STATUS_EARLY:INTEGER);
PORT(A:IN STD_LOGIC_VECTOR(C_WIDTH-1 DOWNTO 0);B:IN STD_LOGIC_VECTOR(C_WIDTH-1 DOWNTO 0):=(OTHERS=>'0');OPERATION:IN
 STD_LOGIC_VECTOR(FLT_PT_OPERATION_WIDTH-1 DOWNTO 0);OPERATION_ND:IN STD_LOGIC;OPERATION_RFD:OUT STD_LOGIC;CLK:IN STD_LOGIC;SCLR:IN
 STD_LOGIC;RESULT:OUT STD_LOGIC_VECTOR(C_WIDTH-1 DOWNTO 0);STATUS:OUT STD_LOGIC_VECTOR(FLT_PT_STATUS_WIDTH-1 DOWNTO 0);EXCEPTION:OUT
 STD_LOGIC;UNDERFLOW:OUT STD_LOGIC;OVERFLOW:OUT STD_LOGIC;INVALID_OP:OUT STD_LOGIC;INEXACT:OUT STD_LOGIC;DIVIDE_BY_ZERO:OUT
 STD_LOGIC;DENORM:OUT STD_LOGIC;RDY:OUT STD_LOGIC);END;ARCHITECTURE BEHAVIORAL OF FLT_PT_OPERATOR IS CONSTANT II1IOOO1II0l1lOl00I1O001I00O0IIIII:INTEGER:=
C_FRACTION_WIDTH;CONSTANT IO1lll0I0l0l1ll1O01Ol0III011IOIIII:INTEGER:=C_WIDTH-C_FRACTION_WIDTH;CONSTANT IOO0111OO0lOOl10l1l000l0OlI0IIIIII:STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII-4 DOWNTO 0):=(OTHERS=>'0');
CONSTANT IIlO1lIIlOlOOO0l10OI1ll0I0O10IIIII:STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0):="10"&IOO0111OO0lOOl10l1l000l0OlI0IIIIII;CONSTANT IOOOlI0llOIl11IO01100OI1llOIIOIIII:STD_LOGIC_VECTOR(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0):=(OTHERS=>'1');
CONSTANT IO1IOOl1111OI1OOII1IOl0lIIIIOIIIII:STD_LOGIC:='1';CONSTANT II1001IO0010Oll1I01lOI0I0IlIOIIIII:STD_LOGIC_VECTOR(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0):=(OTHERS=>'1');CONSTANT IO110I1O0010OIOlIO00l1IIOl0llIIIII:STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII
-2 DOWNTO 0):=(OTHERS=>'0');CONSTANT IIIOOIO01011011IOIIlllIIOO0l1IIIII:STD_LOGIC_VECTOR(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0):=(OTHERS=>'0');CONSTANT II1IOOO00I0OI0O01I000O100llOOIIIII:STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2
 DOWNTO 0):=(OTHERS=>'0');CONSTANT II00OI0110lI1II101lO1OO00I10OIIIII:INTEGER:=2**(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1)-1;CONSTANT II00OIlIlO101I0IIOO0O1I0ll0OIIIIII:INTEGER:=2-2**(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1);CONSTANT IOOI1l1OO01O111lO010OlO1O0l0IIIIII:
INTEGER:=2**(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1)-1;CONSTANT IO11OllII1lO110Ol0I0O00I01l00IIIII:STD_LOGIC_VECTOR:=CONV_STD_LOGIC_VECTOR(2**(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1)-1,IO1lll0I0l0l1ll1O01Ol0III011IOIIII+2);CONSTANT III01lO1l00IOOO0O0I0O0I111O0IIIIII:STD_LOGIC_VECTOR
:=CONV_STD_LOGIC_VECTOR(2**(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1)-1,IO1lll0I0l0l1ll1O01Ol0III011IOIIII+2);CONSTANT IO1I1l01l1OI111Ol0IO10110I11IOIIII:STD_LOGIC_VECTOR:=CONV_STD_LOGIC_VECTOR(2-2**(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1),IO1lll0I0l0l1ll1O01Ol0III011IOIIII+2);PROCEDURE
 IOOll1I1OOlO0lOO0IIII1lO11IIlIIIII(IIIOI11O0OO00OllOllO00lOI000IOIIII:IN INTEGER;IIOIOOO11l0lO001OI10I0IIIIlIIIIIII:IN STD_LOGIC;II0IO0I0Olll01OOO0lIOO01lOlIOOIIII:IN STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0);IOO10IlOOIIIlOIO1IOI1l1lOIIlOIIIII:OUT STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0
);II0l0OlOIIIO1I0IOlIIllOIOO10lIIIII,IO0lIOlI0II1000IOlOIlOI1lIlOOIIIII,IO0O10O101OOIOOl10lIIO101lIIIIIIII:OUT STD_LOGIC)IS VARIABLE IIOl10001I1Ol001OIO01IO1II10OIIIII:STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII DOWNTO 0);VARIABLE IIIO0lOII1OIlOOIO1IlI1lIIO001IIIII:STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1
 DOWNTO 0);VARIABLE IIIIl1100lOI0I1OO1I00OlI0l10IIIIII,IOlI00I100IOOOl011O11IOI1l010IIIII,IIIO1O1110Oll10OI110OIIO111OOIIIII:STD_LOGIC:='0';VARIABLE IIl0OIlO00I0lI101l1I0lO1II0IlIIIII:SIGNED(II1IOOO1II0l1lOl00I1O001I00O0IIIII DOWNTO 0);VARIABLE IOIlII1I0O0l1l1O110O0IOlO0O1lIIIII:INTEGER;VARIABLE
 II11I0011I0IIIl0100l1O01O01O0IIIII:INTEGER;VARIABLE II011lO0O1l10O0I0OIOO000I0O1IOIIII:STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII DOWNTO 0);VARIABLE IO1IIIl1OO00II0ll110l0l0IIO0lIIIII:STD_LOGIC;VARIABLE IIlOllOOI0ll11O1101IIl0l11ll1IIIII:INTEGER;VARIABLE II1I0lOOIIOI1l0l10l0O0l0Ol0OIIIIII:
SIGNED(II1IOOO1II0l1lOl00I1O001I00O0IIIII+3 DOWNTO 0);BEGIN IIIIl1100lOI0I1OO1I00OlI0l10IIIIII:='0';IOlI00I100IOOOl011O11IOI1l010IIIII:='0';IIIO1O1110Oll10OI110OIIO111OOIIIII:='0';II1I0lOOIIOI1l0l10l0O0l0Ol0OIIIIII:=(OTHERS=>'0');IIOl10001I1Ol001OIO01IO1II10OIIIII:=(OTHERS=>'0');II11I0011I0IIIl0100l1O01O01O0IIIII:=CONV_INTEGER(II0IO0I0Olll01OOO0lIOO01lOlIOOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII
+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1)XOR IIOIOOO11l0lO001OI10I0IIIIlIIIIIII);IF IIIOI11O0OO00OllOllO00lOI000IOIIII=1 THEN II11I0011I0IIIl0100l1O01O01O0IIIII:=1-II11I0011I0IIIl0100l1O01O01O0IIIII;END IF;IF II0IO0I0Olll01OOO0lIOO01lOlIOOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1)=IOOOlI0llOIl11IO01100OI1llOIIOIIII AND II0IO0I0Olll01OOO0lIOO01lOlIOOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0)/=IO110I1O0010OIOlIO00l1IIOl0llIIIII THEN
 IIIO0lOII1OIlOOIO1IlI1lIIO001IIIII:=IO1IOOl1111OI1OOII1IOl0lIIIIOIIIII&IOOOlI0llOIl11IO01100OI1llOIIOIIII&IIlO1lIIlOlOOO0l10OI1ll0I0O10IIIII;ELSIF II0IO0I0Olll01OOO0lIOO01lOlIOOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1)=IIIOOIO01011011IOIIlllIIOO0l1IIIII THEN IIIO0lOII1OIlOOIO1IlI1lIIO001IIIII:=CONV_STD_LOGIC_VECTOR(II11I0011I0IIIl0100l1O01O01O0IIIII,1)&IIIOOIO01011011IOIIlllIIOO0l1IIIII&
II1IOOO00I0OI0O01I000O100llOOIIIII;ELSIF II11I0011I0IIIl0100l1O01O01O0IIIII=1 THEN IIIIl1100lOI0I1OO1I00OlI0l10IIIIII:='1';IIIO0lOII1OIlOOIO1IlI1lIIO001IIIII:=IO1IOOl1111OI1OOII1IOl0lIIIIOIIIII&IOOOlI0llOIl11IO01100OI1llOIIOIIII&IIlO1lIIlOlOOO0l10OI1ll0I0O10IIIII;ELSIF II0IO0I0Olll01OOO0lIOO01lOlIOOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1)=II1001IO0010Oll1I01lOI0I0IlIOIIIII AND II0IO0I0Olll01OOO0lIOO01lOlIOOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0
)=IO110I1O0010OIOlIO00l1IIOl0llIIIII THEN IIIO0lOII1OIlOOIO1IlI1lIIO001IIIII:=CONV_STD_LOGIC_VECTOR(II11I0011I0IIIl0100l1O01O01O0IIIII,1)&II1001IO0010Oll1I01lOI0I0IlIOIIIII&IO110I1O0010OIOlIO00l1IIOl0llIIIII;ELSE IIl0OIlO00I0lI101l1I0lO1II0IlIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII):='1';IIl0OIlO00I0lI101l1I0lO1II0IlIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-1 DOWNTO 1):=SIGNED(II0IO0I0Olll01OOO0lIOO01lOlIOOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO
 0));IIl0OIlO00I0lI101l1I0lO1II0IlIIIII(0):='0';IOIlII1I0O0l1l1O110O0IOlO0O1lIIIII:=CONV_INTEGER(UNSIGNED(II0IO0I0Olll01OOO0lIOO01lOlIOOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1)));IF II0IO0I0Olll01OOO0lIOO01lOlIOOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1)=IIIOOIO01011011IOIIlllIIOO0l1IIIII THEN IIl0OIlO00I0lI101l1I0lO1II0IlIIIII:=(OTHERS=>'0'
);END IF;IF II11I0011I0IIIl0100l1O01O01O0IIIII=1 THEN IO1IIIl1OO00II0ll110l0l0IIO0lIIIII:='1';ELSE IO1IIIl1OO00II0ll110l0l0IIO0lIIIII:='0';END IF;IIlOllOOI0ll11O1101IIl0l11ll1IIIII:=(IOIlII1I0O0l1l1O110O0IOlO0O1lIIIII+II00OI0110lI1II101lO1OO00I10OIIIII)/2;IF(IOIlII1I0O0l1l1O110O0IOlO0O1lIIIII MOD 2=1)THEN IIl0OIlO00I0lI101l1I0lO1II0IlIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-1
 DOWNTO 0):=IIl0OIlO00I0lI101l1I0lO1II0IlIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII DOWNTO 1);IIl0OIlO00I0lI101l1I0lO1II0IlIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII):='0';END IF;FOR III1OO10l11110IO1IO0lOII0OO11IIIII IN(II1IOOO1II0l1lOl00I1O001I00O0IIIII)DOWNTO 0 LOOP II1I0lOOIIOI1l0l10l0O0l0Ol0OIIIIII:=II1I0lOOIIOI1l0l10l0O0l0Ol0OIIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+1 DOWNTO 0)&SIGNED(IIl0OIlO00I0lI101l1I0lO1II0IlIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1));IF
 II1I0lOOIIOI1l0l10l0O0l0Ol0OIIIIII>=0 THEN II1I0lOOIIOI1l0l10l0O0l0Ol0OIIIIII:=II1I0lOOIIOI1l0l10l0O0l0Ol0OIIIIII-SIGNED(EXT((IIOl10001I1Ol001OIO01IO1II10OIIIII&"01"),II1IOOO1II0l1lOl00I1O001I00O0IIIII+3));ELSE II1I0lOOIIOI1l0l10l0O0l0Ol0OIIIIII:=II1I0lOOIIOI1l0l10l0O0l0Ol0OIIIIII+SIGNED(EXT((IIOl10001I1Ol001OIO01IO1II10OIIIII&"11"),II1IOOO1II0l1lOl00I1O001I00O0IIIII+3));END IF;IF II1I0lOOIIOI1l0l10l0O0l0Ol0OIIIIII>=0 THEN IIOl10001I1Ol001OIO01IO1II10OIIIII:=IIOl10001I1Ol001OIO01IO1II10OIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-1 DOWNTO 0)&'1';ELSE
 IIOl10001I1Ol001OIO01IO1II10OIIIII:=IIOl10001I1Ol001OIO01IO1II10OIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-1 DOWNTO 0)&'0';END IF;IIl0OIlO00I0lI101l1I0lO1II0IlIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII DOWNTO 0):=IIl0OIlO00I0lI101l1I0lO1II0IlIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0)&"00";END LOOP;IF(IIOl10001I1Ol001OIO01IO1II10OIIIII(0)='1')THEN II011lO0O1l10O0I0OIOO000I0O1IOIIII:=UNSIGNED(EXT(IIOl10001I1Ol001OIO01IO1II10OIIIII
(II1IOOO1II0l1lOl00I1O001I00O0IIIII DOWNTO 1),II1IOOO1II0l1lOl00I1O001I00O0IIIII+1))+1;ELSE II011lO0O1l10O0I0OIOO000I0O1IOIIII:=UNSIGNED(EXT(IIOl10001I1Ol001OIO01IO1II10OIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII DOWNTO 1),II1IOOO1II0l1lOl00I1O001I00O0IIIII+1))+0;END IF;IF(IIlOllOOI0ll11O1101IIl0l11ll1IIIII-II00OI0110lI1II101lO1OO00I10OIIIII)<II00OIlIlO101I0IIOO0O1I0ll0OIIIIII THEN IIIO0lOII1OIlOOIO1IlI1lIIO001IIIII:=
'0'&IIIOOIO01011011IOIIlllIIOO0l1IIIII&II1IOOO00I0OI0O01I000O100llOOIIIII;IIIO1O1110Oll10OI110OIIO111OOIIIII:='1';ELSE IIIO0lOII1OIlOOIO1IlI1lIIO001IIIII:=IO1IIIl1OO00II0ll110l0l0IIO0lIIIII&CONV_STD_LOGIC_VECTOR(IIlOllOOI0ll11O1101IIl0l11ll1IIIII,IO1lll0I0l0l1ll1O01Ol0III011IOIIII)&II011lO0O1l10O0I0OIOO000I0O1IOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0);END IF;END IF
;IOO10IlOOIIIlOIO1IOI1l1lOIIlOIIIII:=IIIO0lOII1OIlOOIO1IlI1lIIO001IIIII;II0l0OlOIIIO1I0IOlIIllOIOO10lIIIII:=IIIIl1100lOI0I1OO1I00OlI0l10IIIIII;IO0lIOlI0II1000IOlOIlOI1lIlOOIIIII:=IOlI00I100IOOOl011O11IOI1l010IIIII;IO0O10O101OOIOOl10lIIO101lIIIIIIII:=IIIO1O1110Oll10OI110OIIO111OOIIIII;END;PROCEDURE IO1O1llOO0IlllI1O1OlOI010l1IIIIIII(IO1O0llO0I1lI11I1O10I0l1O0l0IIIIII:IN INTEGER;II1IO01lI1IO1OII11O1II01I0llIOIIII
:IN INTEGER;II1lIII001001Il0l0OOl0I00I01IIIIII:IN STD_LOGIC;II0O0l0l00OIOl0Ol101Il1Ol0I1lIIIII:IN STD_LOGIC;IOII100I0I1l010IOI1lO1O1I1101IIIII:IN STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0);IOO10OI11Il110I11IIIIIOIO10OlIIIII:IN STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0);IOO1I1lI11Ol1l1OOlllIIII1l1IOIIIII:
OUT STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0);IOl0l10lI11IO10lI1OI1IOI01OO0IIIII,IOO1l1010O10O10I0llO11O100O1IOIIII,IOIlOIOl1lO1l001Ol10IO01OIlI1IIIII,II0IOOI1Il101lO1O010O0O0IO10IOIIII:OUT STD_LOGIC)IS VARIABLE IO1lIIIOl1IIIO1O1lllOO0I1lO0OIIIII,IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII,II111OIOII1IIOOOlO1I011OI0I0lIIIII:
STD_LOGIC_VECTOR(IO1lll0I0l0l1ll1O01Ol0III011IOIIII+1 DOWNTO 0);VARIABLE III0OI0OlIOOl1Ol1I0l00O0lI1IIIIIII,IIIIlI10IO0IlIll11O0O1OII0OIIOIIII,IIIO10O1ll1l0O0IOl0l1lllO0lI1IIIII:STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII-1 DOWNTO 0);VARIABLE IIIlOO0OOl101Ol0Oll10O1lOIIO0IIIII,IIl1O1I0001l1001OllOOII0I10l1IIIII,IIlIlll0III10I0Il0I0OOOIOIIOOIIIII:STD_LOGIC;
VARIABLE IOOI10l0O1lIlIll00Ol1lll10IIIIIIII,IO0OOOI1IIIlIOIIOO0Il00I1lOOlIIIII,IOl0I10010lIIIl000I1O1IO1IlOIIIIII,IOl1I1O0IIO001llOlll1I1lOI1l0IIIII:BOOLEAN;VARIABLE IOl1Ol11IlIl0110l0OOll000lI11IIIII,II001Il0III1O1OI001IOI100000OIIIII,IOOl0llO0OI110111OIOlOIO0lOOIOIIII,II1IOO1l1I11I1ll1OI1I00lII000IIIII:BOOLEAN;CONSTANT II0II1IO1I0IOIl0ll1I0O00lIIOOIIIII:INTEGER:=2;VARIABLE IOOl0IOOO1011llOIOl01lIOI0O11IIIII:STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+
IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0);VARIABLE IIOlOO00Ol0011IIIIIO1I1lllIO0IIIII,II1I0O0100lIIII11lI00l0OOII0lIIIII:STD_LOGIC;VARIABLE IIOIOI0lO1lO100O11Il0OII11OlOIIIII,IO0IlO1lI10Il011101l101IIl0IOIIIII:STD_LOGIC;VARIABLE IOI1O00I10101l0I1001llOOI0I0IOIIII:
STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII-1+II0II1IO1I0IOIl0ll1I0O00lIIOOIIIII+1 DOWNTO 0);VARIABLE IIOIO000I1OI0OlOI1OIOI1l0I0l1IIIII:STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII-1 DOWNTO 0);VARIABLE IO1Il1I0OOOOIl0IOO011l1I0111OIIIII:STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+1 DOWNTO 0);
VARIABLE IO0l0IOllOl1100O10O1O1l0lIO1OIIIII:STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+1 DOWNTO 0);VARIABLE IIlOO000I01110Ill0l1OI1l10IOIOIIII,II1011O1IO1l0llOI11lIIOIlOlIlIIIII,IOO0I1l1IOO0II0O00I0IllOOI1OOIIIII:STD_LOGIC;VARIABLE IOI01l1I0000lIO0IIO01IlIO1001IIIII:STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+1 DOWNTO 0);VARIABLE
 IOI0IIll0I0l1IO0I01lO110IIIIIOIIII:STD_LOGIC;VARIABLE IO00l1I0I1IOlII011Il0l0lOI0OIIIIII:STD_LOGIC;BEGIN IIOlOO00Ol0011IIIIIO1I1lllIO0IIIII:='0';II1I0O0100lIIII11lI00l0OOII0lIIIII:='0';IIOIOI0lO1lO100O11Il0OII11OlOIIIII:='0';IO0IlO1lI10Il011101l101IIl0IOIIIII:='0';IIIlOO0OOl101Ol0Oll10O1lOIIO0IIIII
:=IOII100I0I1l010IOI1lO1O1I1101IIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII+II1IOOO1II0l1lOl00I1O001I00O0IIIII-1);IO1lIIIOl1IIIO1O1lllOO0I1lO0OIIIII:=EXT(IOII100I0I1l010IOI1lO1O1I1101IIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII+II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1),IO1lll0I0l0l1ll1O01Ol0III011IOIIII+2);III0OI0OlIOOl1Ol1I0l00O0lI1IIIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0):=IOII100I0I1l010IOI1lO1O1I1101IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0);III0OI0OlIOOl1Ol1I0l00O0lI1IIIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-1):='1';IIl1O1I0001l1001OllOOII0I10l1IIIII:=IOO10OI11Il110I11IIIIIOIO10OlIIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII+II1IOOO1II0l1lOl00I1O001I00O0IIIII-1);IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII
:=EXT(IOO10OI11Il110I11IIIIIOIO10OlIIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII+II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1),IO1lll0I0l0l1ll1O01Ol0III011IOIIII+2);IIIIlI10IO0IlIll11O0O1OII0OIIOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0):=IOO10OI11Il110I11IIIIIOIO10OlIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0);IIIIlI10IO0IlIll11O0O1OII0OIIOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-1):='1';IF((IO1O0llO0I1lI11I1O10I0l1O0l0IIIIII=1)XOR(II1lIII001001Il0l0OOl0I00I01IIIIII='1'))THEN IIIlOO0OOl101Ol0Oll10O1lOIIO0IIIII
:=NOT IIIlOO0OOl101Ol0Oll10O1lOIIO0IIIII;END IF;IF((II1IO01lI1IO1OII11O1II01I0llIOIIII=1)XOR(II0O0l0l00OIOl0Ol101Il1Ol0I1lIIIII='1'))THEN IIl1O1I0001l1001OllOOII0I10l1IIIII:=NOT IIl1O1I0001l1001OllOOII0I10l1IIIII;END IF;IIlIlll0III10I0Il0I0OOOIOIIOOIIIII:=(IIIlOO0OOl101Ol0Oll10O1lOIIO0IIIII XOR IIl1O1I0001l1001OllOOII0I10l1IIIII);IOOI10l0O1lIlIll00Ol1lll10IIIIIIII:=FALSE;IO0OOOI1IIIlIOIIOO0Il00I1lOOlIIIII:=FALSE;IOl0I10010lIIIl000I1O1IO1IlOIIIIII
:=FALSE;IOl1I1O0IIO001llOlll1I1lOI1l0IIIII:=FALSE;IF IO1lIIIOl1IIIO1O1lllOO0I1lO0OIIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0)=IOOOlI0llOIl11IO01100OI1llOIIOIIII THEN IF III0OI0OlIOOl1Ol1I0l00O0lI1IIIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0)=II1IOOO00I0OI0O01I000O100llOOIIIII THEN IOOI10l0O1lIlIll00Ol1lll10IIIIIIII:=TRUE;ELSE IO0OOOI1IIIlIOIIOO0Il00I1lOOlIIIII:=TRUE;END IF;ELSIF
 IO1lIIIOl1IIIO1O1lllOO0I1lO0OIIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0)=IIIOOIO01011011IOIIlllIIOO0l1IIIII THEN IOl0I10010lIIIl000I1O1IO1IlOIIIIII:=TRUE;ELSE IOl1I1O0IIO001llOlll1I1lOI1l0IIIII:=TRUE;END IF;IOl1Ol11IlIl0110l0OOll000lI11IIIII:=FALSE;II001Il0III1O1OI001IOI100000OIIIII:=FALSE;IOOl0llO0OI110111OIOlOIO0lOOIOIIII:=FALSE;II1IOO1l1I11I1ll1OI1I00lII000IIIII:=FALSE;IF IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1
 DOWNTO 0)=IOOOlI0llOIl11IO01100OI1llOIIOIIII THEN IF IIIIlI10IO0IlIll11O0O1OII0OIIOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0)=II1IOOO00I0OI0O01I000O100llOOIIIII THEN IOl1Ol11IlIl0110l0OOll000lI11IIIII:=TRUE;ELSE II001Il0III1O1OI001IOI100000OIIIII:=TRUE;END IF;ELSIF IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0)=IIIOOIO01011011IOIIlllIIOO0l1IIIII
 THEN IOOl0llO0OI110111OIOlOIO0lOOIOIIII:=TRUE;ELSE II1IOO1l1I11I1ll1OI1I00lII000IIIII:=TRUE;END IF;IF(IO0OOOI1IIIlIOIIOO0Il00I1lOOlIIIII OR II001Il0III1O1OI001IOI100000OIIIII)THEN IOO1I1lI11Ol1l1OOlllIIII1l1IOIIIII:='0'&IOOOlI0llOIl11IO01100OI1llOIIOIIII&IIlO1lIIlOlOOO0l10OI1ll0I0O10IIIII;ELSIF IOOI10l0O1lIlIll00Ol1lll10IIIIIIII THEN IF IOl1Ol11IlIl0110l0OOll000lI11IIIII THEN IOO1I1lI11Ol1l1OOlllIIII1l1IOIIIII:='0'&IOOOlI0llOIl11IO01100OI1llOIIOIIII&
IIlO1lIIlOlOOO0l10OI1ll0I0O10IIIII;IIOlOO00Ol0011IIIIIO1I1lllIO0IIIII:='1';ELSIF IOOl0llO0OI110111OIOlOIO0lOOIOIIII THEN IOO1I1lI11Ol1l1OOlllIIII1l1IOIIIII:=IIlIlll0III10I0Il0I0OOOIOIIOOIIIII&II1001IO0010Oll1I01lOI0I0IlIOIIIII&IO110I1O0010OIOlIO00l1IIOl0llIIIII;ELSE IOO1I1lI11Ol1l1OOlllIIII1l1IOIIIII:=IIlIlll0III10I0Il0I0OOOIOIIOOIIIII&II1001IO0010Oll1I01lOI0I0IlIOIIIII&IO110I1O0010OIOlIO00l1IIOl0llIIIII;END IF;ELSIF IOl0I10010lIIIl000I1O1IO1IlOIIIIII THEN IF IOl1Ol11IlIl0110l0OOll000lI11IIIII
 THEN IOO1I1lI11Ol1l1OOlllIIII1l1IOIIIII:=IIlIlll0III10I0Il0I0OOOIOIIOOIIIII&IIIOOIO01011011IOIIlllIIOO0l1IIIII&II1IOOO00I0OI0O01I000O100llOOIIIII;ELSIF IOOl0llO0OI110111OIOlOIO0lOOIOIIII THEN IOO1I1lI11Ol1l1OOlllIIII1l1IOIIIII:='0'&IOOOlI0llOIl11IO01100OI1llOIIOIIII&IIlO1lIIlOlOOO0l10OI1ll0I0O10IIIII;IIOlOO00Ol0011IIIIIO1I1lllIO0IIIII:='1';ELSE IOO1I1lI11Ol1l1OOlllIIII1l1IOIIIII:=IIlIlll0III10I0Il0I0OOOIOIIOOIIIII&IIIOOIO01011011IOIIlllIIOO0l1IIIII&II1IOOO00I0OI0O01I000O100llOOIIIII;END IF
;ELSE IF IOl1Ol11IlIl0110l0OOll000lI11IIIII THEN IOO1I1lI11Ol1l1OOlllIIII1l1IOIIIII:=IIlIlll0III10I0Il0I0OOOIOIIOOIIIII&IIIOOIO01011011IOIIlllIIOO0l1IIIII&II1IOOO00I0OI0O01I000O100llOOIIIII;ELSIF IOOl0llO0OI110111OIOlOIO0lOOIOIIII THEN IOO1I1lI11Ol1l1OOlllIIII1l1IOIIIII:=IIlIlll0III10I0Il0I0OOOIOIIOOIIIII&II1001IO0010Oll1I01lOI0I0IlIOIIIII&IO110I1O0010OIOlIO00l1IIOl0llIIIII;IO0IlO1lI10Il011101l101IIl0IOIIIII:='1';ELSE II111OIOII1IIOOOlO1I011OI0I0lIIIII:=SIGNED(IO1lIIIOl1IIIO1O1lllOO0I1lO0OIIIII)-
SIGNED(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII);IO1Il1I0OOOOIl0IOO011l1I0111OIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-1 DOWNTO 0):=III0OI0OlIOOl1Ol1I0l00O0lI1IIIIIII;IO1Il1I0OOOOIl0IOO011l1I0111OIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+1 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII):=(OTHERS=>'0');IO0l0IOllOl1100O10O1O1l0lIO1OIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-1 DOWNTO 0):=IIIIlI10IO0IlIll11O0O1OII0OIIOIIII;IO0l0IOllOl1100O10O1O1l0lIO1OIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+1 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII):=(OTHERS=>'0')
;FOR IO01l1ll0IlOll0I00lll11l0OllIIIIII IN II1IOOO1II0l1lOl00I1O001I00O0IIIII+II0II1IO1I0IOIl0ll1I0O00lIIOOIIIII DOWNTO 1 LOOP IF IO1Il1I0OOOOIl0IOO011l1I0111OIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+1)='0'THEN IO1Il1I0OOOOIl0IOO011l1I0111OIIIII:=SIGNED(IO1Il1I0OOOOIl0IOO011l1I0111OIIIII)-SIGNED(IO0l0IOllOl1100O10O1O1l0lIO1OIIIII);IOI1O00I10101l0I1001llOOI0I0IOIIII(IO01l1ll0IlOll0I00lll11l0OllIIIIII):='1';ELSE IO1Il1I0OOOOIl0IOO011l1I0111OIIIII:=SIGNED(IO1Il1I0OOOOIl0IOO011l1I0111OIIIII)+SIGNED(IO0l0IOllOl1100O10O1O1l0lIO1OIIIII);IOI1O00I10101l0I1001llOOI0I0IOIIII(IO01l1ll0IlOll0I00lll11l0OllIIIIII):=
'0';END IF;IO1Il1I0OOOOIl0IOO011l1I0111OIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+1 DOWNTO 1):=IO1Il1I0OOOOIl0IOO011l1I0111OIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII DOWNTO 0);IO1Il1I0OOOOIl0IOO011l1I0111OIIIII(0):='0';END LOOP;IF IO1Il1I0OOOOIl0IOO011l1I0111OIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+1)='0'THEN IO1Il1I0OOOOIl0IOO011l1I0111OIIIII:=SIGNED(IO1Il1I0OOOOIl0IOO011l1I0111OIIIII)-SIGNED(IO0l0IOllOl1100O10O1O1l0lIO1OIIIII);IOI1O00I10101l0I1001llOOI0I0IOIIII(0):='1';
ELSE IO1Il1I0OOOOIl0IOO011l1I0111OIIIII:=SIGNED(IO1Il1I0OOOOIl0IOO011l1I0111OIIIII)+SIGNED(IO0l0IOllOl1100O10O1O1l0lIO1OIIIII);IOI1O00I10101l0I1001llOOI0I0IOIIII(0):='0';END IF;IOI1O00I10101l0I1001llOOI0I0IOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+II0II1IO1I0IOIl0ll1I0O00lIIOOIIIII DOWNTO 1):=IOI1O00I10101l0I1001llOOI0I0IOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-1+II0II1IO1I0IOIl0ll1I0O00lIIOOIIIII DOWNTO 0);IOI1O00I10101l0I1001llOOI0I0IOIIII(0):='1';IIlOO000I01110Ill0l1OI1l10IOIOIIII:=IOI1O00I10101l0I1001llOOI0I0IOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+II0II1IO1I0IOIl0ll1I0O00lIIOOIIIII);IF(IIlOO000I01110Ill0l1OI1l10IOIOIIII=
'1')THEN IIOIO000I1OI0OlOI1OIOI1l0I0l1IIIII:=UNSIGNED(IOI1O00I10101l0I1001llOOI0I0IOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+II0II1IO1I0IOIl0ll1I0O00lIIOOIIIII DOWNTO II0II1IO1I0IOIl0ll1I0O00lIIOOIIIII+1))+UNSIGNED(IOI1O00I10101l0I1001llOOI0I0IOIIII(II0II1IO1I0IOIl0ll1I0O00lIIOOIIIII DOWNTO II0II1IO1I0IOIl0ll1I0O00lIIOOIIIII));IOI0IIll0I0l1IO0I01lO110IIIIIOIIII:=IOI1O00I10101l0I1001llOOI0I0IOIIII(II0II1IO1I0IOIl0ll1I0O00lIIOOIIIII);ELSE II111OIOII1IIOOOlO1I011OI0I0lIIIII:=SIGNED(II111OIOII1IIOOOlO1I011OI0I0lIIIII)-1;IIOIO000I1OI0OlOI1OIOI1l0I0l1IIIII:=UNSIGNED(
IOI1O00I10101l0I1001llOOI0I0IOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+II0II1IO1I0IOIl0ll1I0O00lIIOOIIIII-1 DOWNTO II0II1IO1I0IOIl0ll1I0O00lIIOOIIIII))+UNSIGNED(IOI1O00I10101l0I1001llOOI0I0IOIIII(II0II1IO1I0IOIl0ll1I0O00lIIOOIIIII-1 DOWNTO II0II1IO1I0IOIl0ll1I0O00lIIOOIIIII-1));IOI0IIll0I0l1IO0I01lO110IIIIIOIIII:=IOI1O00I10101l0I1001llOOI0I0IOIIII(II0II1IO1I0IOIl0ll1I0O00lIIOOIIIII-1);END IF;IOI01l1I0000lIO0IIO01IlIO1001IIIII:=SIGNED(IO1Il1I0OOOOIl0IOO011l1I0111OIIIII)+SIGNED(IO0l0IOllOl1100O10O1O1l0lIO1OIIIII)-1;IF SIGNED(IOI01l1I0000lIO0IIO01IlIO1001IIIII)<SIGNED
(CONV_STD_LOGIC_VECTOR(0,II1IOOO1II0l1lOl00I1O001I00O0IIIII+2))AND IOI0IIll0I0l1IO0I01lO110IIIIIOIIII='1'THEN IO00l1I0I1IOlII011Il0l0lOI0OIIIIII:='1';ELSE IO00l1I0I1IOlII011Il0l0lOI0OIIIIII:='0';END IF;IF SIGNED(II111OIOII1IIOOOlO1I011OI0I0lIIIII)>SIGNED(III01lO1l00IOOO0O0I0O0I111O0IIIIII)THEN IOOl0IOOO1011llOIOl01lIOI0O11IIIII
:=IIlIlll0III10I0Il0I0OOOIOIIOOIIIII&II1001IO0010Oll1I01lOI0I0IlIOIIIII&IO110I1O0010OIOlIO00l1IIOl0llIIIII;II1I0O0100lIIII11lI00l0OOII0lIIIII:='1';ELSIF SIGNED(II111OIOII1IIOOOlO1I011OI0I0lIIIII)<SIGNED(IO1I1l01l1OI111Ol0IO10110I11IOIIII)THEN IOOl0IOOO1011llOIOl01lIOI0O11IIIII:=IIlIlll0III10I0Il0I0OOOIOIIOOIIIII&IIIOOIO01011011IOIIlllIIOO0l1IIIII&II1IOOO00I0OI0O01I000O100llOOIIIII;IIOIOI0lO1lO100O11Il0OII11OlOIIIII:='1';
ELSE II111OIOII1IIOOOlO1I011OI0I0lIIIII:=SIGNED(II111OIOII1IIOOOlO1I011OI0I0lIIIII)+SIGNED(IO11OllII1lO110Ol0I0O00I01l00IIIII);IOOl0IOOO1011llOIOl01lIOI0O11IIIII:=IIlIlll0III10I0Il0I0OOOIOIIOOIIIII&II111OIOII1IIOOOlO1I011OI0I0lIIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0)&IIOIO000I1OI0OlOI1OIOI1l0I0l1IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0);END IF;IOO1I1lI11Ol1l1OOlllIIII1l1IOIIIII:=IOOl0IOOO1011llOIOl01lIOI0O11IIIII;END IF;END IF;
IOl0l10lI11IO10lI1OI1IOI01OO0IIIII:=IIOlOO00Ol0011IIIIIO1I1lllIO0IIIII;II0IOOI1Il101lO1O010O0O0IO10IOIIII:=IO0IlO1lI10Il011101l101IIl0IOIIIII;IOO1l1010O10O10I0llO11O100O1IOIIII:=II1I0O0100lIIII11lI00l0OOII0lIIIII;IOIlOIOl1lO1l001Ol10IO01OIlI1IIIII:=IIOIOI0lO1lO100O11Il0OII11OlOIIIII;END;PROCEDURE
 IOI11IOIlOI1II1Il11OlI01Illl0IIIII(IIlO0IOl0I0I0lI0OOll1l1l1lO0IIIIII:IN INTEGER;IOlIOOI0O1OIlOl01O0OIII10O11lIIIII:IN INTEGER;IO1OIOI0I1l11O0IllIOllII1llIIOIIII:IN STD_LOGIC;IIOOO0OOIll110IlI1111I1001I01IIIII:IN STD_LOGIC;IO00lII1lIll0OllOlI1l1O0OI100IIIII:IN STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO
 0);IIII1llIll1l01O1l1O0OIlO1l00OIIIII:IN STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0);II10ll00IlO1IIOIOIO10II0lI1l0IIIII:OUT STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0);IOIIOIIO1lIIOOl0IlO11I00II110IIIII,II0Ol0OI111lIO001O0IIlO110IlIOIIII,II1ll00lO01110lOI1I0IOO0IlO0IIIIII:OUT STD_LOGIC)IS
 VARIABLE IO0I011OOl0OOO000O0I0O0OO0OllIIIII,IO1OllI0IIll0OIOI1l01I010OOIOOIIII,IIOl11l1l101llOl0l0l101I1O1llIIIII:STD_LOGIC_VECTOR(IO1lll0I0l0l1ll1O01Ol0III011IOIIII+1 DOWNTO 0);VARIABLE III1O0Ol0IOOO0IllIOOO000O1lO0IIIII,IIl1IIO111llI0l1O1OI00lIl1I0OIIIII,IIIOOI1II1O11lOIOlOIlOOII1010IIIII:STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII-1 DOWNTO 0);VARIABLE IO0I0I00IO00I1O0I0O0OIOOOI11IOIIII,IIlIOIlO1lO1l1I0OOOI1O1l0O0IOIIIII,IOOI0OO0l1O1O000lO10OOllOIIIIOIIII:STD_LOGIC;
VARIABLE IO1IllOO0II1ll1OII0OOO10OO0I1IIIII:STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+II1IOOO1II0l1lOl00I1O001I00O0IIIII-1 DOWNTO 0);VARIABLE IOOll1I1OO10IlOI0lOO1lOl1O10IOIIII:STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+II1IOOO1II0l1lOl00I1O001I00O0IIIII-1 DOWNTO 0);VARIABLE IOOIOOO1OIO1O0OIIOlOOIOlI1l1lIIIII:STD_LOGIC;VARIABLE
 II10110Oll1OOlIOlOlIl01111IlOIIIII:STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII DOWNTO 0);VARIABLE IOIO00lO11l0IOO1l0I101I11l1OOIIIII:STD_LOGIC_VECTOR(IO1lll0I0l0l1ll1O01Ol0III011IOIIII+1+II1IOOO1II0l1lOl00I1O001I00O0IIIII DOWNTO 0):=(OTHERS=>'0');VARIABLE IIIIl0I1lO1llIOIOOO1lOl11IIlOIIIII:STD_LOGIC_VECTOR(IO1lll0I0l0l1ll1O01Ol0III011IOIIII
+1+II1IOOO1II0l1lOl00I1O001I00O0IIIII DOWNTO 0):=(OTHERS=>'1');VARIABLE II0l0O0IOlIOI00OIl0IlOlI01OI1IIIII,IIlO0l11I10OOIl000I0OOIO0IO0IIIIII:STD_LOGIC;VARIABLE IIOIOOI1ll1O0I1011l0O1lI0IllIOIIII,IOIlllIIlI1OlI0l101llI0II1O1IOIIII:STD_LOGIC;VARIABLE IOO0IO0OOOOO0I10II0llO10ll1OlIIIII,
IIlIII1OIIl0OOl00I0IlOOI1IIlOIIIII:STD_LOGIC;VARIABLE IOl10OI01O100l1IIIl0IIl1lO10lIIIII,IOI1l0OI1IO0llll1llO11Ol1IIlIIIIII:STD_LOGIC;VARIABLE IO00l1II1l000l0I11O010I1IlOlIOIIII,II0IO0O1III0I1I1OlI0011O001IOIIIII:STD_LOGIC;VARIABLE IIl1OOO111O0O11l1OOllOIIIIIl0IIIII,IO00O1llIl1l1I1IIOl11OIlI1lIOOIIII:STD_LOGIC;VARIABLE IOl1I001lIl1Il1I11lI00l11O1OOIIIII,IOlO1OI10Il1OllOl1IIOOIO0I1lIIIIII,III0l0O0I11OOO1lI0OOIO0llOlIlIIIII
:STD_LOGIC;VARIABLE IOO01101I01OlOIO111IIl0OOIOI0IIIII,II00l0IOI1lIlOlOOI0I011O1110OIIIII,IOIO1OI0IlI1I1010lO000IO01Ol0IIIII:STD_LOGIC;VARIABLE IIO00Il10lI0OOllOOO0lO11lOOlIOIIII,IIIIOOlIIO11011I1IlOO10OOOO0OIIIII:STD_LOGIC;BEGIN IO0I011OOl0OOO000O0I0O0OO0OllIIIII:=EXT(IO00lII1lIll0OllOlI1l1O0OI100IIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII+II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1),IO1lll0I0l0l1ll1O01Ol0III011IOIIII+2);IO0I0I00IO00I1O0I0O0OIOOOI11IOIIII:=IO00lII1lIll0OllOlI1l1O0OI100IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII
+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1);III1O0Ol0IOOO0IllIOOO000O1lO0IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0):=IO00lII1lIll0OllOlI1l1O0OI100IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0);III1O0Ol0IOOO0IllIOOO000O1lO0IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-1):='1';IO1OllI0IIll0OIOI1l01I010OOIOOIIII:=EXT(IIII1llIll1l01O1l1O0OIlO1l00OIIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII+II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1),IO1lll0I0l0l1ll1O01Ol0III011IOIIII+2);IIlIOIlO1lO1l1I0OOOI1O1l0O0IOIIIII:=IIII1llIll1l01O1l1O0OIlO1l00OIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1);IIl1IIO111llI0l1O1OI00lIl1I0OIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0):=IIII1llIll1l01O1l1O0OIlO1l00OIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII
-2 DOWNTO 0);IIl1IIO111llI0l1O1OI00lIl1I0OIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-1):='1';IF((IIlO0IOl0I0I0lI0OOll1l1l1lO0IIIIII=1)XOR(IO1OIOI0I1l11O0IllIOllII1llIIOIIII='1'))THEN IO0I0I00IO00I1O0I0O0OIOOOI11IOIIII:=NOT IO0I0I00IO00I1O0I0O0OIOOOI11IOIIII;END IF;IF((IOlIOOI0O1OIlOl01O0OIII10O11lIIIII=1)XOR(IIOOO0OOIll110IlI1111I1001I01IIIII='1'))THEN IIlIOIlO1lO1l1I0OOOI1O1l0O0IOIIIII:=NOT IIlIOIlO1lO1l1I0OOOI1O1l0O0IOIIIII;END IF
;IOOI0OO0l1O1O000lO10OOllOIIIIOIIII:=(IO0I0I00IO00I1O0I0O0OIOOOI11IOIIII XOR IIlIOIlO1lO1l1I0OOOI1O1l0O0IOIIIII);IF IO0I011OOl0OOO000O0I0O0OO0OllIIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0)=IOIO00lO11l0IOO1l0I101I11l1OOIIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0)AND III1O0Ol0IOOO0IllIOOO000O1lO0IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0)=IOIO00lO11l0IOO1l0I101I11l1OOIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0)THEN IIl1OOO111O0O11l1OOllOIIIIIl0IIIII:='1';ELSE IIl1OOO111O0O11l1OOllOIIIIIl0IIIII:='0';
END IF;IF IO1OllI0IIll0OIOI1l01I010OOIOOIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0)=IOIO00lO11l0IOO1l0I101I11l1OOIIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0)AND IIl1IIO111llI0l1O1OI00lIl1I0OIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0)=IOIO00lO11l0IOO1l0I101I11l1OOIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0)THEN IO00O1llIl1l1I1IIOl11OIlI1lIOOIIII:='1';ELSE IO00O1llIl1l1I1IIOl11OIlI1lIOOIIII:='0';END IF;IF III1O0Ol0IOOO0IllIOOO000O1lO0IIIII
(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0)=IOIO00lO11l0IOO1l0I101I11l1OOIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0)THEN II0l0O0IOlIOI00OIl0IlOlI01OI1IIIII:='1';ELSE II0l0O0IOlIOI00OIl0IlOlI01OI1IIIII:='0';END IF;IF IIl1IIO111llI0l1O1OI00lIl1I0OIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0)=IOIO00lO11l0IOO1l0I101I11l1OOIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0)THEN
 IIlO0l11I10OOIl000I0OOIO0IO0IIIIII:='1';ELSE IIlO0l11I10OOIl000I0OOIO0IO0IIIIII:='0';END IF;IF IO0I011OOl0OOO000O0I0O0OO0OllIIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0)=IIIIl0I1lO1llIOIOOO1lOl11IIlOIIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0)THEN IOO0IO0OOOOO0I10II0llO10ll1OlIIIII:='1';ELSE IOO0IO0OOOOO0I10II0llO10ll1OlIIIII:='0';END IF;IF IO1OllI0IIll0OIOI1l01I010OOIOOIIII
(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0)=IIIIl0I1lO1llIOIOOO1lOl11IIlOIIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0)THEN IIlIII1OIIl0OOl00I0IlOOI1IIlOIIIII:='1';ELSE IIlIII1OIIl0OOl00I0IlOOI1IIlOIIIII:='0';END IF;IF IOO0IO0OOOOO0I10II0llO10ll1OlIIIII='1'AND NOT(II0l0O0IOlIOI00OIl0IlOlI01OI1IIIII='1')THEN IOl10OI01O100l1IIIl0IIl1lO10lIIIII:='1';
ELSE IOl10OI01O100l1IIIl0IIl1lO10lIIIII:='0';END IF;IF IIlIII1OIIl0OOl00I0IlOOI1IIlOIIIII='1'AND NOT(IIlO0l11I10OOIl000I0OOIO0IO0IIIIII='1')THEN IOI1l0OI1IO0llll1llO11Ol1IIlIIIIII:='1';ELSE IOI1l0OI1IO0llll1llO11Ol1IIlIIIIII:='0';END IF;IF IOO0IO0OOOOO0I10II0llO10ll1OlIIIII='1'AND II0l0O0IOlIOI00OIl0IlOlI01OI1IIIII='1'THEN
 IO00l1II1l000l0I11O010I1IlOlIOIIII:='1';ELSE IO00l1II1l000l0I11O010I1IlOlIOIIII:='0';END IF;IF IIlIII1OIIl0OOl00I0IlOOI1IIlOIIIII='1'AND IIlO0l11I10OOIl000I0OOIO0IO0IIIIII='1'THEN II0IO0O1III0I1I1OlI0011O001IOIIIII:='1';ELSE II0IO0O1III0I1I1OlI0011O001IOIIIII:='0';END IF;IOIO1OI0IlI1I1010lO000IO01Ol0IIIII:='0';IOO01101I01OlOIO111IIl0OOIOI0IIIII:='0';II00l0IOI1lIlOlOOI0I011O1110OIIIII
:='0';IOl1I001lIl1Il1I11lI00l11O1OOIIIII:='0';IOlO1OI10Il1OllOl1IIOOIO0I1lIIIIII:='0';III0l0O0I11OOO1lI0OOIO0llOlIlIIIII:='0';IF IOl10OI01O100l1IIIl0IIl1lO10lIIIII='1'OR IOI1l0OI1IO0llll1llO11Ol1IIlIIIIII='1'THEN IOl1I001lIl1Il1I11lI00l11O1OOIIIII:='1';ELSIF(IO00l1II1l000l0I11O010I1IlOlIOIIII='1'AND IO00O1llIl1l1I1IIOl11OIlI1lIOOIIII='1')OR(II0IO0O1III0I1I1OlI0011O001IOIIIII='1'AND IIl1OOO111O0O11l1OOllOIIIIIl0IIIII='1')THEN
 IOl1I001lIl1Il1I11lI00l11O1OOIIIII:='1';IOIO1OI0IlI1I1010lO000IO01Ol0IIIII:='1';ELSIF IO00l1II1l000l0I11O010I1IlOlIOIIII='1'OR II0IO0O1III0I1I1OlI0011O001IOIIIII='1'THEN IOlO1OI10Il1OllOl1IIOOIO0I1lIIIIII:='1';ELSIF IIl1OOO111O0O11l1OOllOIIIIIl0IIIII='1'OR IO00O1llIl1l1I1IIOl11OIlI1lIOOIIII='1'THEN III0l0O0I11OOO1lI0OOIO0llOlIlIIIII:='1';ELSE IIOl11l1l101llOl0l0l101I1O1llIIIII:=SIGNED(IO0I011OOl0OOO000O0I0O0OO0OllIIIII)+
SIGNED(IO1OllI0IIll0OIOI1l01I010OOIOOIIII)+1-II00OI0110lI1II101lO1OO00I10OIIIII;IO1IllOO0II1ll1OII0OOO10OO0I1IIIII:=UNSIGNED(III1O0Ol0IOOO0IllIOOO000O1lO0IIIII)*UNSIGNED(IIl1IIO111llI0l1O1OI00lIl1I0OIIIII);IF IO1IllOO0II1ll1OII0OOO10OO0I1IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+II1IOOO1II0l1lOl00I1O001I00O0IIIII-1)='0'THEN IOOll1I1OO10IlOI0lOO1lOl1O10IOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+II1IOOO1II0l1lOl00I1O001I00O0IIIII-1 DOWNTO 0):=IO1IllOO0II1ll1OII0OOO10OO0I1IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0)&'0';IIOl11l1l101llOl0l0l101I1O1llIIIII
:=SIGNED(IIOl11l1l101llOl0l0l101I1O1llIIIII)-1;ELSE IOOll1I1OO10IlOI0lOO1lOl1O10IOIIII:=IO1IllOO0II1ll1OII0OOO10OO0I1IIIII;END IF;IF(IOOll1I1OO10IlOI0lOO1lOl1O10IOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0)=IOIO00lO11l0IOO1l0I101I11l1OOIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0))THEN IOOIOOO1OIO1O0OIIOlOOIOlI1l1lIIIII:='1';ELSE IOOIOOO1OIO1O0OIIOlOOIOlI1l1lIIIII:='0';END IF;IF(IOOll1I1OO10IlOI0lOO1lOl1O10IOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-1)=
'1'AND IOOIOOO1OIO1O0OIIOlOOIOlI1l1lIIIII='0')OR(IOOll1I1OO10IlOI0lOO1lOl1O10IOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-1)='1'AND IOOIOOO1OIO1O0OIIOlOOIOlI1l1lIIIII='1'AND IOOll1I1OO10IlOI0lOO1lOl1O10IOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII)='1')THEN II10110Oll1OOlIOlOlIl01111IlOIIIII:=UNSIGNED(EXT(IOOll1I1OO10IlOI0lOO1lOl1O10IOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+II1IOOO1II0l1lOl00I1O001I00O0IIIII-1 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII),II1IOOO1II0l1lOl00I1O001I00O0IIIII+1))+1;ELSE II10110Oll1OOlIOlOlIl01111IlOIIIII:=EXT
(IOOll1I1OO10IlOI0lOO1lOl1O10IOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+II1IOOO1II0l1lOl00I1O001I00O0IIIII-1 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII),II1IOOO1II0l1lOl00I1O001I00O0IIIII+1);END IF;IF II10110Oll1OOlIOlOlIl01111IlOIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII)='1'THEN IIIOOI1II1O11lOIOlOIlOOII1010IIIII:=II10110Oll1OOlIOlOlIl01111IlOIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII DOWNTO 1);IIOl11l1l101llOl0l0l101I1O1llIIIII:=SIGNED(IIOl11l1l101llOl0l0l101I1O1llIIIII)+1;ELSE IIIOOI1II1O11lOIOlOIlOOII1010IIIII:=II10110Oll1OOlIOlOlIl01111IlOIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-1 DOWNTO 0);END IF;
IOO01101I01OlOIO111IIl0OOIOI0IIIII:='0';II00l0IOI1lIlOlOOI0I011O1110OIIIII:='0';IF SIGNED(IIOl11l1l101llOl0l0l101I1O1llIIIII)<=SIGNED(IOIO00lO11l0IOO1l0I101I11l1OOIIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII+1 DOWNTO 0))THEN III0l0O0I11OOO1lI0OOIO0llOlIlIIIII:='1';II00l0IOI1lIlOlOOI0I011O1110OIIIII:='1';ELSIF IIOl11l1l101llOl0l0l101I1O1llIIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII+1 DOWNTO IO1lll0I0l0l1ll1O01Ol0III011IOIIII)="01"OR(IIOl11l1l101llOl0l0l101I1O1llIIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1
 DOWNTO 0)=NOT IOIO00lO11l0IOO1l0I101I11l1OOIIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0))THEN IOlO1OI10Il1OllOl1IIOOIO0I1lIIIIII:='1';IOO01101I01OlOIO111IIl0OOIOI0IIIII:='1';END IF;END IF;IF IOl1I001lIl1Il1I11lI00l11O1OOIIIII='1'OR IOlO1OI10Il1OllOl1IIOOIO0I1lIIIIII='1'THEN IIOl11l1l101llOl0l0l101I1O1llIIIII:=NOT IOIO00lO11l0IOO1l0I101I11l1OOIIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII+1 DOWNTO 0);IF
 IOl1I001lIl1Il1I11lI00l11O1OOIIIII='1'THEN IIIOOI1II1O11lOIOlOIlOOII1010IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0):=IIlO1lIIlOlOOO0l10OI1ll0I0O10IIIII;ELSE IIIOOI1II1O11lOIOlOIlOOII1010IIIII:=(OTHERS=>'0');END IF;ELSIF III0l0O0I11OOO1lI0OOIO0llOlIlIIIII='1'THEN IIOl11l1l101llOl0l0l101I1O1llIIIII:=(OTHERS=>'0');IIIOOI1II1O11lOIOlOIlOOII1010IIIII:=(OTHERS=>'0');END
 IF;II10ll00IlO1IIOIOIO10II0lI1l0IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0):=IOOI0OO0l1O1O000lO10OOllOIIIIOIIII&IIOl11l1l101llOl0l0l101I1O1llIIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0)&IIIOOI1II1O11lOIOlOIlOOII1010IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0);II0Ol0OI111lIO001O0IIlO110IlIOIIII:=IOO01101I01OlOIO111IIl0OOIOI0IIIII;II1ll00lO01110lOI1I0IOO0IlO0IIIIII:=II00l0IOI1lIlOlOOI0I011O1110OIIIII;IOIIOIIO1lIIOOl0IlO11I00II110IIIII:=IOIO1OI0IlI1I1010lO000IO01Ol0IIIII;END;PROCEDURE
 IIO0101IlI11I0IOlI01l1ll0O10OIIIII(IOl00OIO0IOOllO1I1O101lIIl11OIIIII:IN INTEGER;IOl011Ol0O1Il1IIIIlIOlIl101IlIIIII:IN INTEGER;IO00OI0ll1l1l0llI1I000OOO0010IIIII:IN STD_LOGIC;IOl0OIIOl0O00OO0lI0I0O1IO1OOIOIIII:IN STD_LOGIC;IOI0111Il0IllIIO0O0lO0I111010IIIII:IN STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0);IOO0IOIOOll0Il0OlI001lIIIOOOIIIIII
:IN STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0);IOO0llOIlIO0110l1lOO01I00l1OIIIIII:OUT STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0);IOIO0OOIOIOl0OIllO011O11O0OOIIIIII,IO0lI0OlO11O10O1III000O01l0l0IIIII,IIO1O00llO01OII1I11lIIO001lI0IIIII:OUT STD_LOGIC)IS
 CONSTANT IOIl1lI1IO111IO0OII101O1I0l0IOIIII:SIGNED(II1IOOO1II0l1lOl00I1O001I00O0IIIII-1 DOWNTO 0):=(OTHERS=>'0');CONSTANT IOOIOOOlO000O1I0lOI1OO01l0OOlIIIII:SIGNED(II1IOOO1II0l1lOl00I1O001I00O0IIIII DOWNTO 0):='1'&IOIl1lI1IO111IO0OII101O1I0l0IOIIII;CONSTANT
 IO01O100lOO0IOOI000OO1lIOO1l0IIIII:SIGNED(II1IOOO1II0l1lOl00I1O001I00O0IIIII DOWNTO 0):=(OTHERS=>'0');CONSTANT IOl1100I00OlIllOI1I0III1O1l01IIIII:SIGNED(II1IOOO1II0l1lOl00I1O001I00O0IIIII DOWNTO 0):=(OTHERS=>'0');CONSTANT IO1OlIO1l10Ill0O11IO0I0ll1OlIIIIII:SIGNED(2
*II1IOOO1II0l1lOl00I1O001I00O0IIIII+3-1 DOWNTO 0):=IO01O100lOO0IOOI000OO1lIOO1l0IIIII&'1'&IOl1100I00OlIllOI1I0III1O1l01IIIII;CONSTANT IIOIlOO1lI01O10O1Ol0OOI10110OIIIII:SIGNED(2*II1IOOO1II0l1lOl00I1O001I00O0IIIII+2 DOWNTO 0):=(OTHERS=>'0');VARIABLE IO0II1lll1llOlO1lll1001O1IlOIOIIII:
STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0);VARIABLE IOOO00lOlO0l0llI01lIlOOIIllIlIIIII,IIlIIII1lOllO0IlO11I1O01110IOIIIII,II0I1I1l00l1O11OOIOIIllII10IlIIIII:STD_LOGIC;VARIABLE III0lIIOOIOl0ll0ll0l1lO10IlIIIIIII:SIGNED(2*II1IOOO1II0l1lOl00I1O001I00O0IIIII+2 DOWNTO 0);VARIABLE
 III010I1Ol1OlOI0IO10O0000II11IIIII:SIGNED(2*II1IOOO1II0l1lOl00I1O001I00O0IIIII+2 DOWNTO 0);VARIABLE IOIlOO00I1I00lO00l0I00OlIO01IIIIII:INTEGER;VARIABLE IIO111Il00001lO0l00lOOlI1IO10IIIII:INTEGER;VARIABLE II10IOlI11OOI1IO1OlI0IlI0I0I1IIIII:INTEGER;VARIABLE IO1lO1OOOl00OOI0lOI1Ol1O1lI0IIIIII:INTEGER;
VARIABLE IO0I10OO0llIIlII1I01OOI001IIIIIIII:INTEGER;VARIABLE II110IlI0l101IO1IlI1O00llI00OIIIII:SIGNED(2*II1IOOO1II0l1lOl00I1O001I00O0IIIII+2 DOWNTO 0);VARIABLE III0O000IO1IOIO10l0I00lOIII11IIIII:STD_LOGIC;VARIABLE II1llIOlOlll00O010O1lI1IOI1I1IIIII:INTEGER;VARIABLE
 IO1I11OIllI1III1III11OlIIlIIOIIIII:INTEGER;BEGIN IOOO00lOlO0l0llI01lIlOOIIllIlIIIII:='0';IIlIIII1lOllO0IlO11I1O01110IOIIIII:='0';II0I1I1l00l1O11OOIOIIllII10IlIIIII:='0';IO1lO1OOOl00OOI0lOI1Ol1O1lI0IIIIII:=CONV_INTEGER(IOI0111Il0IllIIO0O0lO0I111010IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1)XOR IO00OI0ll1l1l0llI1I000OOO0010IIIII);IF IOl00OIO0IOOllO1I1O101lIIl11OIIIII=1 THEN
 IO1lO1OOOl00OOI0lOI1Ol1O1lI0IIIIII:=1-IO1lO1OOOl00OOI0lOI1Ol1O1lI0IIIIII;END IF;IO0I10OO0llIIlII1I01OOI001IIIIIIII:=CONV_INTEGER(IOO0IOIOOll0Il0OlI001lIIIOOOIIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1)XOR IOl0OIIOl0O00OO0lI0I0O1IO1OOIOIIII);IF IOl011Ol0O1Il1IIIIlIOlIl101IlIIIII=1 THEN IO0I10OO0llIIlII1I01OOI001IIIIIIII:=1-IO0I10OO0llIIlII1I01OOI001IIIIIIII;END IF;IF IOI0111Il0IllIIO0O0lO0I111010IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1)=
IIIOOIO01011011IOIIlllIIOO0l1IIIII AND IOO0IOIOOll0Il0OlI001lIIIOOOIIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1)=IIIOOIO01011011IOIIlllIIOO0l1IIIII THEN IF(IO1lO1OOOl00OOI0lOI1Ol1O1lI0IIIIII+IO0I10OO0llIIlII1I01OOI001IIIIIIII)=2 THEN III0O000IO1IOIO10l0I00lOIII11IIIII:='1';ELSE III0O000IO1IOIO10l0I00lOIII11IIIII:='0';END IF;IO0II1lll1llOlO1lll1001O1IlOIOIIII:=III0O000IO1IOIO10l0I00lOIII11IIIII&
IIIOOIO01011011IOIIlllIIOO0l1IIIII&II1IOOO00I0OI0O01I000O100llOOIIIII;ELSIF IOI0111Il0IllIIO0O0lO0I111010IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1)=IOOOlI0llOIl11IO01100OI1llOIIOIIII AND IOI0111Il0IllIIO0O0lO0I111010IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0)/=IO110I1O0010OIOlIO00l1IIOl0llIIIII THEN IO0II1lll1llOlO1lll1001O1IlOIOIIII:=IO1IOOl1111OI1OOII1IOl0lIIIIOIIIII&IOOOlI0llOIl11IO01100OI1llOIIOIIII&IIlO1lIIlOlOOO0l10OI1ll0I0O10IIIII;ELSIF IOO0IOIOOll0Il0OlI001lIIIOOOIIIIII(
II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1)=IOOOlI0llOIl11IO01100OI1llOIIOIIII AND IOO0IOIOOll0Il0OlI001lIIIOOOIIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0)/=IO110I1O0010OIOlIO00l1IIOl0llIIIII THEN IO0II1lll1llOlO1lll1001O1IlOIOIIII:=IO1IOOl1111OI1OOII1IOl0lIIIIOIIIII&IOOOlI0llOIl11IO01100OI1llOIIOIIII&IIlO1lIIlOlOOO0l10OI1ll0I0O10IIIII;ELSIF IOI0111Il0IllIIO0O0lO0I111010IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1)=
II1001IO0010Oll1I01lOI0I0IlIOIIIII AND IOI0111Il0IllIIO0O0lO0I111010IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0)=IO110I1O0010OIOlIO00l1IIOl0llIIIII AND IOO0IOIOOll0Il0OlI001lIIIOOOIIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1)=II1001IO0010Oll1I01lOI0I0IlIOIIIII AND IOO0IOIOOll0Il0OlI001lIIIOOOIIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0)=IO110I1O0010OIOlIO00l1IIOl0llIIIII THEN IF IO1lO1OOOl00OOI0lOI1Ol1O1lI0IIIIII=IO0I10OO0llIIlII1I01OOI001IIIIIIII THEN IO0II1lll1llOlO1lll1001O1IlOIOIIII
:=CONV_STD_LOGIC_VECTOR(IO1lO1OOOl00OOI0lOI1Ol1O1lI0IIIIII,1)&II1001IO0010Oll1I01lOI0I0IlIOIIIII&IO110I1O0010OIOlIO00l1IIOl0llIIIII;ELSE IO0II1lll1llOlO1lll1001O1IlOIOIIII:=IO1IOOl1111OI1OOII1IOl0lIIIIOIIIII&IOOOlI0llOIl11IO01100OI1llOIIOIIII&IIlO1lIIlOlOOO0l10OI1ll0I0O10IIIII;IOOO00lOlO0l0llI01lIlOOIIllIlIIIII:='1';END IF;ELSIF IOI0111Il0IllIIO0O0lO0I111010IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-2 DOWNTO
 II1IOOO1II0l1lOl00I1O001I00O0IIIII-1)=II1001IO0010Oll1I01lOI0I0IlIOIIIII AND IOI0111Il0IllIIO0O0lO0I111010IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0)=IO110I1O0010OIOlIO00l1IIOl0llIIIII THEN IO0II1lll1llOlO1lll1001O1IlOIOIIII:=CONV_STD_LOGIC_VECTOR(IO1lO1OOOl00OOI0lOI1Ol1O1lI0IIIIII,1)&II1001IO0010Oll1I01lOI0I0IlIOIIIII&IO110I1O0010OIOlIO00l1IIOl0llIIIII;ELSIF IOO0IOIOOll0Il0OlI001lIIIOOOIIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1
)=II1001IO0010Oll1I01lOI0I0IlIOIIIII AND IOO0IOIOOll0Il0OlI001lIIIOOOIIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0)=IO110I1O0010OIOlIO00l1IIOl0llIIIII THEN IO0II1lll1llOlO1lll1001O1IlOIOIIII:=CONV_STD_LOGIC_VECTOR(IO0I10OO0llIIlII1I01OOI001IIIIIIII,1)&II1001IO0010Oll1I01lOI0I0IlIOIIIII&IO110I1O0010OIOlIO00l1IIOl0llIIIII;ELSE III0lIIOOIOl0ll0ll0l1lO10IlIIIIIII:=(OTHERS=>'0');III0lIIOOIOl0ll0ll0l1lO10IlIIIIIII(2
*II1IOOO1II0l1lOl00I1O001I00O0IIIII):='1';III0lIIOOIOl0ll0ll0l1lO10IlIIIIIII(2*II1IOOO1II0l1lOl00I1O001I00O0IIIII-1 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII+1):=SIGNED(IOI0111Il0IllIIO0O0lO0I111010IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0));IOIlOO00I1I00lO00l0I00OlIO01IIIIII:=CONV_INTEGER(UNSIGNED(IOI0111Il0IllIIO0O0lO0I111010IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1)));IOIlOO00I1I00lO00l0I00OlIO01IIIIII:=IOIlOO00I1I00lO00l0I00OlIO01IIIIII-
II00OI0110lI1II101lO1OO00I10OIIIII;III010I1Ol1OlOI0IO10O0000II11IIIII:=(OTHERS=>'0');III010I1Ol1OlOI0IO10O0000II11IIIII(2*II1IOOO1II0l1lOl00I1O001I00O0IIIII):='1';III010I1Ol1OlOI0IO10O0000II11IIIII(2*II1IOOO1II0l1lOl00I1O001I00O0IIIII-1 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII+1):=SIGNED(IOO0IOIOOll0Il0OlI001lIIIOOOIIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0));IIO111Il00001lO0l00lOOlI1IO10IIIII:=CONV_INTEGER(UNSIGNED(IOO0IOIOOll0Il0OlI001lIIIOOOIIIIII
(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1)));IIO111Il00001lO0l00lOOlI1IO10IIIII:=IIO111Il00001lO0l00lOOlI1IO10IIIII-II00OI0110lI1II101lO1OO00I10OIIIII;IF IOI0111Il0IllIIO0O0lO0I111010IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1)=IIIOOIO01011011IOIIlllIIOO0l1IIIII THEN III0lIIOOIOl0ll0ll0l1lO10IlIIIIIII:=(OTHERS=>'0');END IF;IF IOO0IOIOOll0Il0OlI001lIIIOOOIIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-2
 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1)=IIIOOIO01011011IOIIlllIIOO0l1IIIII THEN III010I1Ol1OlOI0IO10O0000II11IIIII:=(OTHERS=>'0');END IF;IF IOIlOO00I1I00lO00l0I00OlIO01IIIIII>IIO111Il00001lO0l00lOOlI1IO10IIIII THEN II10IOlI11OOI1IO1OlI0IlI0I0I1IIIII:=IOIlOO00I1I00lO00l0I00OlIO01IIIIII-IIO111Il00001lO0l00lOOlI1IO10IIIII;II1llIOlOlll00O010O1lI1IOI1I1IIIII:=IOIlOO00I1I00lO00l0I00OlIO01IIIIII;III010I1Ol1OlOI0IO10O0000II11IIIII:=SHR(III010I1Ol1OlOI0IO10O0000II11IIIII,
CONV_UNSIGNED(II10IOlI11OOI1IO1OlI0IlI0I0I1IIIII,IO1lll0I0l0l1ll1O01Ol0III011IOIIII+1));ELSE II10IOlI11OOI1IO1OlI0IlI0I0I1IIIII:=IIO111Il00001lO0l00lOOlI1IO10IIIII-IOIlOO00I1I00lO00l0I00OlIO01IIIIII;II1llIOlOlll00O010O1lI1IOI1I1IIIII:=IIO111Il00001lO0l00lOOlI1IO10IIIII;III0lIIOOIOl0ll0ll0l1lO10IlIIIIIII:=SHR(III0lIIOOIOl0ll0ll0l1lO10IlIIIIIII,CONV_UNSIGNED(II10IOlI11OOI1IO1OlI0IlI0I0I1IIIII,IO1lll0I0l0l1ll1O01Ol0III011IOIIII+1));END IF;IF
 IO1lO1OOOl00OOI0lOI1Ol1O1lI0IIIIII=0 THEN IF IO0I10OO0llIIlII1I01OOI001IIIIIIII=0 THEN II110IlI0l101IO1IlI1O00llI00OIIIII:=III0lIIOOIOl0ll0ll0l1lO10IlIIIIIII+III010I1Ol1OlOI0IO10O0000II11IIIII;ELSE II110IlI0l101IO1IlI1O00llI00OIIIII:=III0lIIOOIOl0ll0ll0l1lO10IlIIIIIII-III010I1Ol1OlOI0IO10O0000II11IIIII;END IF;ELSE IF IO0I10OO0llIIlII1I01OOI001IIIIIIII=0 THEN II110IlI0l101IO1IlI1O00llI00OIIIII:=III010I1Ol1OlOI0IO10O0000II11IIIII-III0lIIOOIOl0ll0ll0l1lO10IlIIIIIII;ELSE
 II110IlI0l101IO1IlI1O00llI00OIIIII:=-(III0lIIOOIOl0ll0ll0l1lO10IlIIIIIII+III010I1Ol1OlOI0IO10O0000II11IIIII);END IF;END IF;IF II110IlI0l101IO1IlI1O00llI00OIIIII(2*II1IOOO1II0l1lOl00I1O001I00O0IIIII+2)='1'THEN II110IlI0l101IO1IlI1O00llI00OIIIII:=ABS(II110IlI0l101IO1IlI1O00llI00OIIIII);III0O000IO1IOIO10l0I00lOIII11IIIII:='1';ELSE III0O000IO1IOIO10l0I00lOIII11IIIII:='0';END IF;IF
 II110IlI0l101IO1IlI1O00llI00OIIIII(2*II1IOOO1II0l1lOl00I1O001I00O0IIIII+1)='1'THEN II110IlI0l101IO1IlI1O00llI00OIIIII:=SHR(II110IlI0l101IO1IlI1O00llI00OIIIII,CONV_UNSIGNED(1,1));II1llIOlOlll00O010O1lI1IOI1I1IIIII:=II1llIOlOlll00O010O1lI1IOI1I1IIIII+1;ELSE IO1I11OIllI1III1III11OlIIlIIOIIIII:=0;WHILE IO1I11OIllI1III1III11OlIIlIIOIIIII<2*II1IOOO1II0l1lOl00I1O001I00O0IIIII AND
 II110IlI0l101IO1IlI1O00llI00OIIIII(2*II1IOOO1II0l1lOl00I1O001I00O0IIIII)='0'LOOP II110IlI0l101IO1IlI1O00llI00OIIIII:=SHL(II110IlI0l101IO1IlI1O00llI00OIIIII,CONV_UNSIGNED(1,1));IO1I11OIllI1III1III11OlIIlIIOIIIII:=IO1I11OIllI1III1III11OlIIlIIOIIIII+1;END LOOP;II1llIOlOlll00O010O1lI1IOI1I1IIIII:=II1llIOlOlll00O010O1lI1IOI1I1IIIII-IO1I11OIllI1III1III11OlIIlIIOIIIII;END IF
;IF II110IlI0l101IO1IlI1O00llI00OIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII)='0'THEN ELSIF II110IlI0l101IO1IlI1O00llI00OIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII DOWNTO 0)=IOOIOOOlO000O1I0lOI1OO01l0OOlIIIII THEN IF II110IlI0l101IO1IlI1O00llI00OIIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII+1)='1'THEN II110IlI0l101IO1IlI1O00llI00OIIIII:=II110IlI0l101IO1IlI1O00llI00OIIIII+IO1OlIO1l10Ill0O11IO0I0ll1OlIIIIII;ELSE END IF;
ELSE II110IlI0l101IO1IlI1O00llI00OIIIII:=II110IlI0l101IO1IlI1O00llI00OIIIII+IO1OlIO1l10Ill0O11IO0I0ll1OlIIIIII;END IF;IF II110IlI0l101IO1IlI1O00llI00OIIIII(2*II1IOOO1II0l1lOl00I1O001I00O0IIIII+1)='1'THEN II110IlI0l101IO1IlI1O00llI00OIIIII:=SHR(II110IlI0l101IO1IlI1O00llI00OIIIII,CONV_UNSIGNED(1,1));II1llIOlOlll00O010O1lI1IOI1I1IIIII:=II1llIOlOlll00O010O1lI1IOI1I1IIIII+1;END IF
;IF II110IlI0l101IO1IlI1O00llI00OIIIII=IIOIlOO1lI01O10O1Ol0OOI10110OIIIII THEN IO0II1lll1llOlO1lll1001O1IlOIOIIII:='0'&IIIOOIO01011011IOIIlllIIOO0l1IIIII&II1IOOO00I0OI0O01I000O100llOOIIIII;ELSIF II1llIOlOlll00O010O1lI1IOI1I1IIIII<II00OIlIlO101I0IIOO0O1I0ll0OIIIIII THEN IO0II1lll1llOlO1lll1001O1IlOIOIIII:=III0O000IO1IOIO10l0I00lOIII11IIIII&IIIOOIO01011011IOIIlllIIOO0l1IIIII&II1IOOO00I0OI0O01I000O100llOOIIIII;II0I1I1l00l1O11OOIOIIllII10IlIIIII:='1'
;ELSIF II1llIOlOlll00O010O1lI1IOI1I1IIIII>IOOI1l1OO01O111lO010OlO1O0l0IIIIII THEN IO0II1lll1llOlO1lll1001O1IlOIOIIII:=III0O000IO1IOIO10l0I00lOIII11IIIII&II1001IO0010Oll1I01lOI0I0IlIOIIIII&IO110I1O0010OIOlIO00l1IIOl0llIIIII;IIlIIII1lOllO0IlO11I1O01110IOIIIII:='1';ELSE II1llIOlOlll00O010O1lI1IOI1I1IIIII:=II1llIOlOlll00O010O1lI1IOI1I1IIIII+II00OI0110lI1II101lO1OO00I10OIIIII;IO0II1lll1llOlO1lll1001O1IlOIOIIII:=III0O000IO1IOIO10l0I00lOIII11IIIII&
CONV_STD_LOGIC_VECTOR(II1llIOlOlll00O010O1lI1IOI1I1IIIII,IO1lll0I0l0l1ll1O01Ol0III011IOIIII)&CONV_STD_LOGIC_VECTOR(II110IlI0l101IO1IlI1O00llI00OIIIII(2*II1IOOO1II0l1lOl00I1O001I00O0IIIII-1 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII+1),II1IOOO1II0l1lOl00I1O001I00O0IIIII-1);END IF;END IF;IOO0llOIlIO0110l1lOO01I00l1OIIIIII:=IO0II1lll1llOlO1lll1001O1IlOIOIIII;IOIO0OOIOIOl0OIllO011O11O0OOIIIIII:=
IOOO00lOlO0l0llI01lIlOOIIllIlIIIII;IO0lI0OlO11O10O1III000O01l0l0IIIII:=IIlIIII1lOllO0IlO11I1O01110IOIIIII;IIO1O00llO01OII1I11lIIO001lI0IIIII:=II0I1I1l00l1O11OOIOIIllII10IlIIIII;END;PROCEDURE IIl11lIlOO0IIII0IOlI0l1000I1IIIIII(IOOI10l11llO01llIIllOI1IO0l1OIIIII:IN INTEGER;IOO1IIll11IlI110IOlllI1Il1IO1IIIII:IN INTEGER;IOO000O0Ol1OlIOOI00l11I1l1I00IIIII:IN
 STD_LOGIC;IIll0O11l1O1lOl111IIOlOIl0I0OIIIII:IN STD_LOGIC;IIOI10lI0II00O0IOOl0I10001lO1IIIII:IN STD_LOGIC_VECTOR(FLT_PT_COMPARE_OPERATION_WIDTH-1 DOWNTO 0);IIO1IIOOO0OO1100OO11l0OOllIIIOIIII:IN STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1
 DOWNTO 0);IOO01O011lIIIlOl1O0lOIOOI110IOIIII:IN STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0);IOIOO101OO01Ol1101l1O01O1OOllIIIII:OUT STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0);IIOO0IIlO0O0I01l00I1011II0011IIIII:OUT STD_LOGIC)IS VARIABLE
 IOl0lOIIO0IllIOIO1Oll0lOOOII1IIIII:UNSIGNED(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0);VARIABLE IIOlI0O00IO011lIIOl100O001lIOOIIII:UNSIGNED(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0);VARIABLE III0IlIOll1Ill0I0I0OlIO10I1I1IIIII:UNSIGNED(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0);VARIABLE IOOllIl0I1ll0lII0IOIIO1lI10IIIIIII:UNSIGNED
(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0);VARIABLE II0I1O11OOll0l0I11O110OlI0lIOOIIII:STD_LOGIC;VARIABLE II1lI1l0l00llI0l0l1O0OOII10I1IIIII:STD_LOGIC;VARIABLE II0l10llII1lO0O1lOIlOOI10I0lIIIIII:BOOLEAN;VARIABLE IO1I1OlOI1OII110llI1lI0IIl0O0IIIII:BOOLEAN;VARIABLE II110IO0lllI1lOI110IO00I1lOlIIIIII:
BOOLEAN;VARIABLE IIl110lllO10l0llOI11l01I0I1OlIIIII:BOOLEAN;VARIABLE IOOll11IO1O1llOIl10010O1IIOOIIIIII:STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0);VARIABLE IIII00I101O111lII1O000IO1lOOIIIIII:BOOLEAN;VARIABLE
 IOOI01II11O1I1IOII1II01O1001lIIIII:BOOLEAN;VARIABLE IO111Il1I1O0lO1OlOI0l01I1O010IIIII:STD_LOGIC;BEGIN II0I1O11OOll0l0I11O110OlI0lIOOIIII:=IIO1IIOOO0OO1100OO11l0OOllIIIOIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII+II1IOOO1II0l1lOl00I1O001I00O0IIIII-1);III0IlIOll1Ill0I0I0OlIO10I1I1IIIII:=UNSIGNED(IIO1IIOOO0OO1100OO11l0OOllIIIOIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII+II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1));IOl0lOIIO0IllIOIO1Oll0lOOOII1IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO
 0):=UNSIGNED(IIO1IIOOO0OO1100OO11l0OOllIIIOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0));II1lI1l0l00llI0l0l1O0OOII10I1IIIII:=IOO01O011lIIIlOl1O0lOIOOI110IOIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII+II1IOOO1II0l1lOl00I1O001I00O0IIIII-1);IOOllIl0I1ll0lII0IOIIO1lI10IIIIIII:=UNSIGNED(IOO01O011lIIIlOl1O0lOIOOI110IOIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII+II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1));IIOlI0O00IO011lIIOl100O001lIOOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0):=UNSIGNED(IOO01O011lIIIlOl1O0lOIOOI110IOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2
 DOWNTO 0));IF((IOOI10l11llO01llIIllOI1IO0l1OIIIII=1)XOR(IOO000O0Ol1OlIOOI00l11I1l1I00IIIII='1'))THEN II0I1O11OOll0l0I11O110OlI0lIOOIIII:=NOT II0I1O11OOll0l0I11O110OlI0lIOOIIII;END IF;IF((IOO1IIll11IlI110IOlllI1Il1IO1IIIII=1)XOR(IIll0O11l1O1lOl111IIOlOIl0I0OIIIII='1'))THEN II1lI1l0l00llI0l0l1O0OOII10I1IIIII:=NOT II1lI1l0l00llI0l0l1O0OOII10I1IIIII;END IF;
II0l10llII1lO0O1lOIlOOI10I0lIIIIII:=FALSE;IO1I1OlOI1OII110llI1lI0IIl0O0IIIII:=FALSE;II110IO0lllI1lOI110IO00I1lOlIIIIII:=FALSE;IIl110lllO10l0llOI11l01I0I1OlIIIII:=FALSE;IO111Il1I1O0lO1OlOI0l01I1O010IIIII:='0';IF(II0I1O11OOll0l0I11O110OlI0lIOOIIII='0'AND II1lI1l0l00llI0l0l1O0OOII10I1IIIII='1')THEN II110IO0lllI1lOI110IO00I1lOlIIIIII:=TRUE;ELSIF(II0I1O11OOll0l0I11O110OlI0lIOOIIII='1'
AND II1lI1l0l00llI0l0l1O0OOII10I1IIIII='0')THEN IO1I1OlOI1OII110llI1lI0IIl0O0IIIII:=TRUE;ELSIF(III0IlIOll1Ill0I0I0OlIO10I1I1IIIII/=IOOllIl0I1ll0lII0IOIIO1lI10IIIIIII)THEN IF(IOOllIl0I1ll0lII0IOIIO1lI10IIIIIII>III0IlIOll1Ill0I0I0OlIO10I1I1IIIII)THEN IO1I1OlOI1OII110llI1lI0IIl0O0IIIII:=(II0I1O11OOll0l0I11O110OlI0lIOOIIII='0');II110IO0lllI1lOI110IO00I1lOlIIIIII:=(II0I1O11OOll0l0I11O110OlI0lIOOIIII='1');ELSE IO1I1OlOI1OII110llI1lI0IIl0O0IIIII:=(
II0I1O11OOll0l0I11O110OlI0lIOOIIII='1');II110IO0lllI1lOI110IO00I1lOlIIIIII:=(II0I1O11OOll0l0I11O110OlI0lIOOIIII='0');END IF;ELSE IF(IIOlI0O00IO011lIIOl100O001lIOOIIII>IOl0lOIIO0IllIOIO1Oll0lOOOII1IIIII)THEN IO1I1OlOI1OII110llI1lI0IIl0O0IIIII:=(II0I1O11OOll0l0I11O110OlI0lIOOIIII='0');II110IO0lllI1lOI110IO00I1lOlIIIIII:=(II0I1O11OOll0l0I11O110OlI0lIOOIIII='1');ELSE IF(IIOlI0O00IO011lIIOl100O001lIOOIIII/=IOl0lOIIO0IllIOIO1Oll0lOOOII1IIIII)THEN
 IO1I1OlOI1OII110llI1lI0IIl0O0IIIII:=(II0I1O11OOll0l0I11O110OlI0lIOOIIII='1');II110IO0lllI1lOI110IO00I1lOlIIIIII:=(II0I1O11OOll0l0I11O110OlI0lIOOIIII='0');ELSE II0l10llII1lO0O1lOIlOOI10I0lIIIIII:=TRUE;END IF;END IF;END IF;IF(((III0IlIOll1Ill0I0I0OlIO10I1I1IIIII=UNSIGNED(IIIOOIO01011011IOIIlllIIOO0l1IIIII))AND(IOl0lOIIO0IllIOIO1Oll0lOOOII1IIIII=UNSIGNED(
II1IOOO00I0OI0O01I000O100llOOIIIII)))AND((IOOllIl0I1ll0lII0IOIIO1lI10IIIIIII=UNSIGNED(IIIOOIO01011011IOIIlllIIOO0l1IIIII))AND(IIOlI0O00IO011lIIOl100O001lIOOIIII=UNSIGNED(II1IOOO00I0OI0O01I000O100llOOIIIII))))THEN II0l10llII1lO0O1lOIlOOI10I0lIIIIII:=TRUE;IO1I1OlOI1OII110llI1lI0IIl0O0IIIII:=FALSE;II110IO0lllI1lOI110IO00I1lOlIIIIII:=FALSE;END IF;IF(((
III0IlIOll1Ill0I0I0OlIO10I1I1IIIII=UNSIGNED(IOOOlI0llOIl11IO01100OI1llOIIOIIII))AND(IOl0lOIIO0IllIOIO1Oll0lOOOII1IIIII/=UNSIGNED(II1IOOO00I0OI0O01I000O100llOOIIIII)))OR((IOOllIl0I1ll0lII0IOIIO1lI10IIIIIII=UNSIGNED(IOOOlI0llOIl11IO01100OI1llOIIOIIII))AND(IIOlI0O00IO011lIIOl100O001lIOOIIII/=UNSIGNED(II1IOOO00I0OI0O01I000O100llOOIIIII))))THEN II0l10llII1lO0O1lOIlOOI10I0lIIIIII:=
FALSE;IO1I1OlOI1OII110llI1lI0IIl0O0IIIII:=FALSE;II110IO0lllI1lOI110IO00I1lOlIIIIII:=FALSE;IIl110lllO10l0llOI11l01I0I1OlIIIII:=TRUE;END IF;IOOll11IO1O1llOIl10010O1IIOOIIIIII:=(OTHERS=>'0');IF((II110IO0lllI1lOI110IO00I1lOlIIIIII AND(IIOI10lI0II00O0IOOl0I10001lO1IIIII(2)='1'))OR(II0l10llII1lO0O1lOIlOOI10I0lIIIIII AND(IIOI10lI0II00O0IOOl0I10001lO1IIIII(1)=
'1'))OR(IO1I1OlOI1OII110llI1lI0IIl0O0IIIII AND(IIOI10lI0II00O0IOOl0I10001lO1IIIII(0)='1')))THEN IOOll11IO1O1llOIl10010O1IIOOIIIIII(0):='1';END IF;IF(IIOI10lI0II00O0IOOl0I10001lO1IIIII="000")THEN IF(IIl110lllO10l0llOI11l01I0I1OlIIIII)THEN IOOll11IO1O1llOIl10010O1IIOOIIIIII(0):='1';END IF;END IF;IF(((
III0IlIOll1Ill0I0I0OlIO10I1I1IIIII=UNSIGNED(IIIOOIO01011011IOIIlllIIOO0l1IIIII))AND(IOl0lOIIO0IllIOIO1Oll0lOOOII1IIIII/=UNSIGNED(II1IOOO00I0OI0O01I000O100llOOIIIII)))OR((IOOllIl0I1ll0lII0IOIIO1lI10IIIIIII=UNSIGNED(IIIOOIO01011011IOIIlllIIOO0l1IIIII))AND(IIOlI0O00IO011lIIOl100O001lIOOIIII/=UNSIGNED(II1IOOO00I0OI0O01I000O100llOOIIIII))))THEN IOOll11IO1O1llOIl10010O1IIOOIIIIII(0)
:='0';ELSE IIII00I101O111lII1O000IO1lOOIIIIII:=((III0IlIOll1Ill0I0I0OlIO10I1I1IIIII=UNSIGNED(IOOOlI0llOIl11IO01100OI1llOIIOIIII))AND(IOl0lOIIO0IllIOIO1Oll0lOOOII1IIIII/=UNSIGNED(II1IOOO00I0OI0O01I000O100llOOIIIII)))AND(IOl0lOIIO0IllIOIO1Oll0lOOOII1IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2)='0');IOOI01II11O1I1IOII1II01O1001lIIIII:=((IOOllIl0I1ll0lII0IOIIO1lI10IIIIIII=
UNSIGNED(IOOOlI0llOIl11IO01100OI1llOIIOIIII))AND(IIOlI0O00IO011lIIOl100O001lIOOIIII/=UNSIGNED(II1IOOO00I0OI0O01I000O100llOOIIIII)))AND(IIOlI0O00IO011lIIOl100O001lIOOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2)='0');IF((IIII00I101O111lII1O000IO1lOOIIIIII OR IOOI01II11O1I1IOII1II01O1001lIIIII)OR(IIl110lllO10l0llOI11l01I0I1OlIIIII AND NOT(IIOI10lI0II00O0IOOl0I10001lO1IIIII=
"000"OR IIOI10lI0II00O0IOOl0I10001lO1IIIII="010"OR IIOI10lI0II00O0IOOl0I10001lO1IIIII="101")))THEN IO111Il1I1O0lO1OlOI0l01I1O010IIIII:='1';IOOll11IO1O1llOIl10010O1IIOOIIIIII(0):='0';END IF;END IF;IOIOO101OO01Ol1101l1O01O1OOllIIIII:=IOOll11IO1O1llOIl10010O1IIOOIIIIII;IIOO0IIlO0O0I01l00I1011II0011IIIII:=IO111Il1I1O0lO1OlOI0l01I1O010IIIII;END;SIGNAL
 III011IIIl1IO1l0O11000I0llI00IIIII:INTEGER:=2;TYPE II1O1ll0lOO0Ol1O0OO01I0OI0lIIOIIII IS ARRAY(NATURAL RANGE<>)OF STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0);TYPE IIO1l1Ol1l11Il0000II00lI011I0IIIII IS ARRAY(NATURAL RANGE<>)OF
 STD_LOGIC_VECTOR(FLT_PT_OPERATION_WIDTH-1 DOWNTO 0);SIGNAL IIO1OllIOO1lI1OOO1IOIII1lIl0IOIIII:STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0):=(OTHERS=>'0');SIGNAL II1lI11lI1II1000lOllIOl01l0l0IIIII:
STD_LOGIC_VECTOR(II1IOOO1II0l1lOl00I1O001I00O0IIIII+IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0):=(OTHERS=>'0');SIGNAL II0l0001lI0I0IlllI1I100OO10IIIIIII:STD_LOGIC_VECTOR(FLT_PT_OPERATION_WIDTH-1 DOWNTO 0):=(OTHERS
=>'0');CONSTANT II01l0llO10l10II111lIlOIllO0lIIIII:INTEGER:=100;SIGNAL IOl0I1O0OllIl0lI1IlO0OIlII0lIIIIII:II1O1ll0lOO0Ol1O0OO01I0OI0lIIOIIII(0 TO II01l0llO10l10II111lIlOIllO0lIIIII-1);SIGNAL IIlI1l00I0IOl1l1O0llllO0I1I0IIIIII:II1O1ll0lOO0Ol1O0OO01I0OI0lIIOIIII(0 TO
 II01l0llO10l10II111lIlOIllO0lIIIII-1);SIGNAL IIl1O01ll1111l0llIOO0OOl1ll0IOIIII:IIO1l1Ol1l11Il0000II00lI011I0IIIII(0 TO II01l0llO10l10II111lIlOIllO0lIIIII-1);SIGNAL II10l111IOllO0O1111Ill001lll1IIIII:STD_LOGIC_VECTOR(0 TO
 II01l0llO10l10II111lIlOIllO0lIIIII-1):=(OTHERS=>'0');SIGNAL IIlOI1II1OOlOl00Ol01IOl0OO0OOIIIII:STD_LOGIC:='0';SIGNAL IIll1lO0l0lI0OII00l00OO11IlO1IIIII:STD_LOGIC:='0';SIGNAL III00O11l11IlIOI1llIIIOII100lIIIII:
STD_LOGIC:='0';SIGNAL IO1l01O110OIl00l10lOOlI0lI0I0IIIII:STD_LOGIC;SIGNAL IIlIO1lIl0lI1lOlI0I0O0I0OO0IIIIIII:STD_LOGIC:='0';SIGNAL IOIIOO1001lI01IOOlOllIOOIO1O1IIIII:STD_LOGIC;SIGNAL
 IIOlIO1l10OOO1l1IlII1ll0100IOIIIII:STD_LOGIC;SIGNAL III1I01Ill1l0lOIlO01lO0I1IlIIOIIII:STD_LOGIC;SIGNAL IOOIl1OOO1IIl11O00lI1IlOIIl0OIIIII:STD_LOGIC;SIGNAL IOlI00ll1I0I1ll0ll01l1OOl0IlIIIIII:STD_LOGIC;BEGIN
 IO1l01O110OIl00l10lOOlI0lI0I0IIIII<=III00O11l11IlIOI1llIIIOII100lIIIII AND OPERATION_ND AND NOT(SCLR);RDF_CNTRL:PROCESS(CLK)BEGIN IF RISING_EDGE(CLK)THEN IF SCLR='1'THEN
 IIlOI1II1OOlOl00Ol01IOl0OO0OOIIIII<='0';ELSE IIlOI1II1OOlOl00Ol01IOl0OO0OOIIIII<=IIll1lO0l0lI0OII00l00OO11IlO1IIIII;END IF;IF SCLR='1'THEN III00O11l11IlIOI1llIIIOII100lIIIII<='0';IIlIO1lIl0lI1lOlI0I0O0I0OO0IIIIIII<='0';ELSIF
 IIlIO1lIl0lI1lOlI0I0O0I0OO0IIIIIII='1'THEN IF IIll1lO0l0lI0OII00l00OO11IlO1IIIII='1'THEN III00O11l11IlIOI1llIIIOII100lIIIII<='1';IIlIO1lIl0lI1lOlI0I0O0I0OO0IIIIIII<='0';END IF;ELSIF IO1l01O110OIl00l10lOOlI0lI0I0IIIII='1'THEN
 IF((OPERATION(FLT_PT_OP_CODE_SLICE)=FLT_PT_DIVIDE_OP_CODE_SLV)AND(C_OPTIMIZATION=FLT_PT_UNOPTIMIZED))THEN IIlIO1lIl0lI1lOlI0I0O0I0OO0IIIIIII<='1';
III00O11l11IlIOI1llIIIOII100lIIIII<='0';ELSE III00O11l11IlIOI1llIIIOII100lIIIII<='1';END IF;ELSE III00O11l11IlIOI1llIIIOII100lIIIII<='1';END IF;END IF;END PROCESS;III011IIIl1IO1l0O11000I0llI00IIIII<=FLT_PT_DELAY
(FAMILY=>C_FAMILY,OP_CODE=>OPERATION(FLT_PT_OP_CODE_SLICE),WIDTH=>C_WIDTH,FRACTION_WIDTH=>C_FRACTION_WIDTH,OPTIMIZATION=>
C_OPTIMIZATION,MULT_USAGE=>C_MULT_USAGE,RATE=>-1);PROCESS(CLK)BEGIN IF RISING_EDGE(CLK)THEN IF SCLR='1'THEN IOl0I1O0OllIl0lI1IlO0OIlII0lIIIIII<=(OTHERS=>(
OTHERS=>'0'));IIlI1l00I0IOl1l1O0llllO0I1I0IIIIII<=(OTHERS=>(OTHERS=>'0'));IIl1O01ll1111l0llIOO0OOl1ll0IOIIII<=(OTHERS=>(OTHERS=>'0'));ELSE IOl0I1O0OllIl0lI1IlO0OIlII0lIIIIII(0 TO III011IIIl1IO1l0O11000I0llI00IIIII-1)<=A&IOl0I1O0OllIl0lI1IlO0OIlII0lIIIIII(0 TO
 III011IIIl1IO1l0O11000I0llI00IIIII-2);IIlI1l00I0IOl1l1O0llllO0I1I0IIIIII(0 TO III011IIIl1IO1l0O11000I0llI00IIIII-1)<=B&IIlI1l00I0IOl1l1O0llllO0I1I0IIIIII(0 TO III011IIIl1IO1l0O11000I0llI00IIIII-2);IIl1O01ll1111l0llIOO0OOl1ll0IOIIII(0 TO III011IIIl1IO1l0O11000I0llI00IIIII-1)<=OPERATION&IIl1O01ll1111l0llIOO0OOl1ll0IOIIII(0 TO III011IIIl1IO1l0O11000I0llI00IIIII-2);END
 IF;II10l111IOllO0O1111Ill001lll1IIIII(0 TO III011IIIl1IO1l0O11000I0llI00IIIII-1)<=IO1l01O110OIl00l10lOOlI0lI0I0IIIII&II10l111IOllO0O1111Ill001lll1IIIII(0 TO III011IIIl1IO1l0O11000I0llI00IIIII-2);END IF;END PROCESS;IIO1OllIOO1lI1OOO1IOIII1lIl0IOIIII<=IOl0I1O0OllIl0lI1IlO0OIlII0lIIIIII(III011IIIl1IO1l0O11000I0llI00IIIII-1);II1lI11lI1II1000lOllIOl01l0l0IIIII<=IIlI1l00I0IOl1l1O0llllO0I1I0IIIIII(III011IIIl1IO1l0O11000I0llI00IIIII-1
);II0l0001lI0I0IlllI1I100OO10IIIIIII<=IIl1O01ll1111l0llIOO0OOl1ll0IOIIII(III011IIIl1IO1l0O11000I0llI00IIIII-1);IIll1lO0l0lI0OII00l00OO11IlO1IIIII<=II10l111IOllO0O1111Ill001lll1IIIII(III011IIIl1IO1l0O11000I0llI00IIIII-2);PROCESS(IIO1OllIOO1lI1OOO1IOIII1lIl0IOIIII,II1lI11lI1II1000lOllIOl01l0l0IIIII,II0l0001lI0I0IlllI1I100OO10IIIIIII)VARIABLE III11I01Ol11IOO00IOI1I11OOl10IIIII:
STD_LOGIC_VECTOR(C_WIDTH-1 DOWNTO 0);VARIABLE IIl1lOIllIlIl01ll00O11OIl100IOIIII:STD_LOGIC;VARIABLE IIOII0OO1Ol0lOOlO1O1OOlllIllOIIIII:STD_LOGIC;VARIABLE II1011l1lI11IlIlI0l0l00100lO0IIIII:
STD_LOGIC;VARIABLE IO1OO10IOIO11O10IOOOllllI1Il0IIIII:STD_LOGIC;VARIABLE II1IOl1011OlI0O00l1O10OlllOI0IIIII:STD_LOGIC;VARIABLE IO1OIOllI1llI01O00IIl0O111IIOOIIII:BOOLEAN;VARIABLE IO01001lO000lI1lI0IO11lO0I1OlIIIII:BOOLEAN;
VARIABLE IOOl11OIOl101I1I1I00lIlIlO00IIIIII:BOOLEAN;VARIABLE IIlOOO01III1O0O0IOII0I0lOlIlOIIIII:BOOLEAN;VARIABLE IIIl1IO0lOOOIIlOOllOl010IOl1IOIIII:BOOLEAN;VARIABLE IIl010l00OlI0lO1OO11Il10lIOIOOIIII:BOOLEAN;VARIABLE
 IIOIl1I10OOOllIlIOl11lI0IO1lIOIIII:BOOLEAN;BEGIN IIl1lOIllIlIl01ll00O11OIl100IOIIII:='0';IIOII0OO1Ol0lOOlO1O1OOlllIllOIIIII:='0';II1011l1lI11IlIlI0l0l00100lO0IIIII:='0';IO1OO10IOIO11O10IOOOllllI1Il0IIIII:='0';II1IOl1011OlI0O00l1O10OlllOI0IIIII:='0';IIOIl1I10OOOllIlIOl11lI0IO1lIOIIII:=(
FLT_PT_NUMBER_OF_INPUTS(CONV_INTEGER(UNSIGNED(OPERATION(FLT_PT_OP_CODE_SLICE))))=2);IO1OIOllI1llI01O00IIl0O111IIOOIIII:=((IIO1OllIOO1lI1OOO1IOIII1lIl0IOIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII+II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1)=IOOOlI0llOIl11IO01100OI1llOIIOIIII)
AND(IIO1OllIOO1lI1OOO1IOIII1lIl0IOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0)/=II1IOOO00I0OI0O01I000O100llOOIIIII));IO01001lO000lI1lI0IO11lO0I1OlIIIII:=((II1lI11lI1II1000lOllIOl01l0l0IIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII+II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1)=IOOOlI0llOIl11IO01100OI1llOIIOIIII)AND(II1lI11lI1II1000lOllIOl01l0l0IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0)/=II1IOOO00I0OI0O01I000O100llOOIIIII));
IOOl11OIOl101I1I1I00lIlIlO00IIIIII:=IO1OIOllI1llI01O00IIl0O111IIOOIIII AND(IIO1OllIOO1lI1OOO1IOIII1lIl0IOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2)='0');IIlOOO01III1O0O0IOII0I0lOlIlOIIIII:=IO01001lO000lI1lI0IO11lO0I1OlIIIII AND(II1lI11lI1II1000lOllIOl01l0l0IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2)='0');IIIl1IO0lOOOIIlOOllOl010IOl1IOIIII:=((IIO1OllIOO1lI1OOO1IOIII1lIl0IOIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII+II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1)=
IIIOOIO01011011IOIIlllIIOO0l1IIIII)AND(IIO1OllIOO1lI1OOO1IOIII1lIl0IOIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0)/=II1IOOO00I0OI0O01I000O100llOOIIIII));IIl010l00OlI0lO1OO11Il10lIOIOOIIII:=((II1lI11lI1II1000lOllIOl01l0l0IIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII+II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO II1IOOO1II0l1lOl00I1O001I00O0IIIII-1)=IIIOOIO01011011IOIIlllIIOO0l1IIIII)AND(II1lI11lI1II1000lOllIOl01l0l0IIIII(II1IOOO1II0l1lOl00I1O001I00O0IIIII-2 DOWNTO 0)/=II1IOOO00I0OI0O01I000O100llOOIIIII
));IF(IO1OIOllI1llI01O00IIl0O111IIOOIIII OR(IO01001lO000lI1lI0IO11lO0I1OlIIIII AND IIOIl1I10OOOllIlIOl11lI0IO1lIOIIII))THEN III11I01Ol11IOO00IOI1I11OOl10IIIII:=IO1IOOl1111OI1OOII1IOl0lIIIIOIIIII&IOOOlI0llOIl11IO01100OI1llOIIOIIII&IIlO1lIIlOlOOO0l10OI1ll0I0O10IIIII;IIl1lOIllIlIl01ll00O11OIl100IOIIII:='1';IF NOT(IOOl11OIOl101I1I1I00lIlIlO00IIIIII OR(
IIlOOO01III1O0O0IOII0I0lOlIlOIIIII AND IIOIl1I10OOOllIlIOl11lI0IO1lIOIIII))THEN IIl1lOIllIlIl01ll00O11OIl100IOIIII:='0';END IF;ELSIF(IIIl1IO0lOOOIIlOOllOl010IOl1IOIIII OR(IIl010l00OlI0lO1OO11Il10lIOIOOIIII AND IIOIl1I10OOOllIlIOl11lI0IO1lIOIIII))THEN III11I01Ol11IOO00IOI1I11OOl10IIIII:=IO1IOOl1111OI1OOII1IOl0lIIIIOIIIII&
IOOOlI0llOIl11IO01100OI1llOIIOIIII&IIlO1lIIlOlOOO0l10OI1ll0I0O10IIIII;II1IOl1011OlI0O00l1O10OlllOI0IIIII:='1';ELSE CASE CONV_INTEGER(UNSIGNED(II0l0001lI0I0IlllI1I100OO10IIIIIII(FLT_PT_OP_CODE_SLICE)))IS WHEN FLT_PT_SQRT_OP_CODE=>
IOOll1I1OOlO0lOO0IIII1lO11IIlIIIII(0,'0',IIO1OllIOO1lI1OOO1IOIII1lIl0IOIIII,III11I01Ol11IOO00IOI1I11OOl10IIIII,IIl1lOIllIlIl01ll00O11OIl100IOIIII,IIOII0OO1Ol0lOOlO1O1OOlllIllOIIIII,IO1OO10IOIO11O10IOOOllllI1Il0IIIII);WHEN FLT_PT_DIVIDE_OP_CODE=>IO1O1llOO0IlllI1O1OlOI010l1IIIIIII(0,0,'0','0',
IIO1OllIOO1lI1OOO1IOIII1lIl0IOIIII,II1lI11lI1II1000lOllIOl01l0l0IIIII,III11I01Ol11IOO00IOI1I11OOl10IIIII,IIl1lOIllIlIl01ll00O11OIl100IOIIII,IIOII0OO1Ol0lOOlO1O1OOlllIllOIIIII,IO1OO10IOIO11O10IOOOllllI1Il0IIIII,II1011l1lI11IlIlI0l0l00100lO0IIIII);WHEN FLT_PT_MULTIPLY_OP_CODE=>IOI11IOIlOI1II1Il11OlI01Illl0IIIII(0
,0,'0','0',IIO1OllIOO1lI1OOO1IOIII1lIl0IOIIII,II1lI11lI1II1000lOllIOl01l0l0IIIII,III11I01Ol11IOO00IOI1I11OOl10IIIII,IIl1lOIllIlIl01ll00O11OIl100IOIIII,IIOII0OO1Ol0lOOlO1O1OOlllIllOIIIII,IO1OO10IOIO11O10IOOOllllI1Il0IIIII);WHEN FLT_PT_ADD_OP_CODE=>IIO0101IlI11I0IOlI01l1ll0O10OIIIII(0,0,'0','0',IIO1OllIOO1lI1OOO1IOIII1lIl0IOIIII,
II1lI11lI1II1000lOllIOl01l0l0IIIII,III11I01Ol11IOO00IOI1I11OOl10IIIII,IIl1lOIllIlIl01ll00O11OIl100IOIIII,IIOII0OO1Ol0lOOlO1O1OOlllIllOIIIII,IO1OO10IOIO11O10IOOOllllI1Il0IIIII);WHEN FLT_PT_SUBTRACT_OP_CODE=>IIO0101IlI11I0IOlI01l1ll0O10OIIIII(0,0,'0','1',IIO1OllIOO1lI1OOO1IOIII1lIl0IOIIII,II1lI11lI1II1000lOllIOl01l0l0IIIII,
III11I01Ol11IOO00IOI1I11OOl10IIIII,IIl1lOIllIlIl01ll00O11OIl100IOIIII,IIOII0OO1Ol0lOOlO1O1OOlllIllOIIIII,IO1OO10IOIO11O10IOOOllllI1Il0IIIII);WHEN FLT_PT_COMPARE_OP_CODE=>IIl11lIlOO0IIII0IOlI0l1000I1IIIIII(0,0,'0','0',II0l0001lI0I0IlllI1I100OO10IIIIIII(
FLT_PT_COMPARE_OPERATION_SLICE),IIO1OllIOO1lI1OOO1IOIII1lIl0IOIIII,II1lI11lI1II1000lOllIOl01l0l0IIIII,III11I01Ol11IOO00IOI1I11OOl10IIIII,IIl1lOIllIlIl01ll00O11OIl100IOIIII);WHEN OTHERS=>ASSERT(FALSE)REPORT
"Internal error: flt_pt_operation(behavioral)"&" - contact Xilinx support"SEVERITY FAILURE;END CASE;END IF;RESULT<=III11I01Ol11IOO00IOI1I11OOl10IIIII;
IOIIOO1001lI01IOOlOllIOOIO1O1IIIII<=IIl1lOIllIlIl01ll00O11OIl100IOIIII;IIOlIO1l10OOO1l1IlII1ll0100IOIIIII<=IIOII0OO1Ol0lOOlO1O1OOlllIllOIIIII;III1I01Ill1l0lOIlO01lO0I1IlIIOIIII<=IO1OO10IOIO11O10IOOOllllI1Il0IIIII;IOOIl1OOO1IIl11O00lI1IlOIIl0OIIIII<=II1011l1lI11IlIlI0l0l00100lO0IIIII;
IOlI00ll1I0I1ll0ll01l1OOl0IlIIIIII<=II1IOl1011OlI0O00l1O10OlllOI0IIIII;END PROCESS;OPERATION_RFD<=III00O11l11IlIOI1llIIIOII100lIIIII;YES_EARLY:IF C_STATUS_EARLY=FLT_PT_YES GENERATE RDY<=
IIll1lO0l0lI0OII00l00OO11IlO1IIIII;END GENERATE;NO_EARLY:IF C_STATUS_EARLY=FLT_PT_NO GENERATE RDY<=IIlOI1II1OOlOl00Ol01IOl0OO0OOIIIII;END GENERATE;INVALID_OP<=IOIIOO1001lI01IOOlOllIOOIO1O1IIIII;
OVERFLOW<=IIOlIO1l10OOO1l1IlII1ll0100IOIIIII;UNDERFLOW<=III1I01Ill1l0lOIlO01lO0I1IlIIOIIII;DIVIDE_BY_ZERO<=IOOIl1OOO1IIl11O00lI1IlOIIl0OIIIII;DENORM<=IOlI00ll1I0I1ll0ll01l1OOl0IlIIIIII;STATUS<=IOIIOO1001lI01IOOlOllIOOIO1O1IIIII&
IOOIl1OOO1IIl11O00lI1IlOIIl0OIIIII&IIOlIO1l10OOO1l1IlII1ll0100IOIIIII&III1I01Ill1l0lOIlO01lO0I1IlIIOIIII&IOlI00ll1I0I1ll0ll01l1OOl0IlIIIIII;END;LIBRARY IEEE;USE IEEE.STD_LOGIC_1164.ALL;USE IEEE.NUMERIC_STD.ALL;
LIBRARY XILINXCORELIB;USE XILINXCORELIB.FLOATING_POINT_V1_0_CONSTS.ALL;USE XILINXCORELIB.FLOATING_POINT_PKG_V1_0.ALL;ENTITY
 FLOATING_POINT_V1_0_XST IS GENERIC(C_FAMILY:STRING:=C_FAMILY_DEFAULT;C_HAS_ADD:INTEGER:=C_HAS_ADD_DEFAULT;C_HAS_SUBTRACT:INTEGER:=
C_HAS_SUBTRACT_DEFAULT;C_HAS_MULTIPLY:INTEGER:=C_HAS_MULTIPLY_DEFAULT;C_HAS_DIVIDE:INTEGER:=C_HAS_DIVIDE_DEFAULT;C_HAS_SQRT:INTEGER
:=C_HAS_SQRT_DEFAULT;C_HAS_COMPARE:INTEGER:=C_HAS_COMPARE_DEFAULT;C_HAS_FIX_TO_FLT:INTEGER:=C_HAS_FIX_TO_FLT_DEFAULT;
C_HAS_FLT_TO_FIX:INTEGER:=C_HAS_FLT_TO_FIX_DEFAULT;C_A_WIDTH:INTEGER:=C_A_WIDTH_DEFAULT;C_A_FRACTION_WIDTH:INTEGER:=
C_A_FRACTION_WIDTH_DEFAULT;C_B_WIDTH:INTEGER:=C_B_WIDTH_DEFAULT;C_B_FRACTION_WIDTH:INTEGER:=C_B_FRACTION_WIDTH_DEFAULT;
C_RESULT_WIDTH:INTEGER:=C_RESULT_WIDTH_DEFAULT;C_RESULT_FRACTION_WIDTH:INTEGER:=C_RESULT_FRACTION_WIDTH_DEFAULT;C_COMPARE_OPERATION
:INTEGER:=C_COMPARE_OPERATION_DEFAULT;C_LATENCY:INTEGER:=C_LATENCY_DEFAULT;C_OPTIMIZATION:INTEGER:=C_OPTIMIZATION_DEFAULT;
C_MULT_USAGE:INTEGER:=C_MULT_USAGE_DEFAULT;C_RATE:INTEGER:=C_RATE_DEFAULT;C_HAS_ACLR:INTEGER:=C_HAS_ACLR_DEFAULT;C_HAS_CE:INTEGER:=
C_HAS_CE_DEFAULT;C_HAS_SCLR:INTEGER:=C_HAS_SCLR_DEFAULT;C_HAS_A_NEGATE:INTEGER:=C_HAS_A_NEGATE_DEFAULT;C_HAS_B_NEGATE:INTEGER:=
C_HAS_B_NEGATE_DEFAULT;C_HAS_A_ND:INTEGER:=C_HAS_A_ND_DEFAULT;C_HAS_A_RFD:INTEGER:=C_HAS_A_RFD_DEFAULT;C_HAS_B_ND:INTEGER:=
C_HAS_B_ND_DEFAULT;C_HAS_B_RFD:INTEGER:=C_HAS_B_RFD_DEFAULT;C_HAS_OPERATION_ND:INTEGER:=C_HAS_OPERATION_ND_DEFAULT;
C_HAS_OPERATION_RFD:INTEGER:=C_HAS_OPERATION_RFD_DEFAULT;C_HAS_RDY:INTEGER:=C_HAS_RDY_DEFAULT;C_HAS_CTS:INTEGER:=C_HAS_CTS_DEFAULT;
C_HAS_UNDERFLOW:INTEGER:=C_HAS_UNDERFLOW_DEFAULT;C_HAS_OVERFLOW:INTEGER:=C_HAS_OVERFLOW_DEFAULT;C_HAS_INVALID_OP:INTEGER:=
C_HAS_INVALID_OP_DEFAULT;C_HAS_INEXACT:INTEGER:=C_HAS_INEXACT_DEFAULT;C_HAS_DIVIDE_BY_ZERO:INTEGER:=C_HAS_DIVIDE_BY_ZERO_DEFAULT;
C_HAS_STATUS:INTEGER:=C_HAS_STATUS_DEFAULT;C_HAS_EXCEPTION:INTEGER:=C_HAS_EXCEPTION_DEFAULT;C_STATUS_EARLY:INTEGER:=
C_STATUS_EARLY_DEFAULT);PORT(A:IN STD_LOGIC_VECTOR(C_A_WIDTH-1 DOWNTO 0);B:IN STD_LOGIC_VECTOR(C_B_WIDTH-1 DOWNTO 0):=(OTHERS=>'0');
A_NEGATE:IN STD_LOGIC:='0';B_NEGATE:IN STD_LOGIC:='0';OPERATION:IN STD_LOGIC_VECTOR(FLT_PT_OPERATION_WIDTH-1 DOWNTO 0):=(OTHERS=>'0'
);A_ND:IN STD_LOGIC:='1';A_RFD:OUT STD_LOGIC;B_ND:IN STD_LOGIC:='1';B_RFD:OUT STD_LOGIC;OPERATION_ND:IN STD_LOGIC:='1';OPERATION_RFD
:OUT STD_LOGIC;CLK:IN STD_LOGIC;SCLR:IN STD_LOGIC:='0';ACLR:IN STD_LOGIC:='0';CE:IN STD_LOGIC:='1';RESULT:OUT STD_LOGIC_VECTOR(
C_RESULT_WIDTH-1 DOWNTO 0);STATUS:OUT STD_LOGIC_VECTOR(FLT_PT_STATUS_WIDTH-1 DOWNTO 0);EXCEPTION:OUT STD_LOGIC;UNDERFLOW:OUT
 STD_LOGIC;OVERFLOW:OUT STD_LOGIC;INVALID_OP:OUT STD_LOGIC;INEXACT:OUT STD_LOGIC;DIVIDE_BY_ZERO:OUT STD_LOGIC;RDY:OUT STD_LOGIC;CTS
:IN STD_LOGIC:='1');END;ARCHITECTURE BEHAVIORAL OF FLOATING_POINT_V1_0_XST IS COMPONENT FLT_PT_OPERATOR GENERIC(C_FAMILY:STRING;
C_WIDTH:INTEGER;C_FRACTION_WIDTH:INTEGER;C_OPTIMIZATION:INTEGER;C_MULT_USAGE:INTEGER;C_HAS_STATUS:INTEGER;C_STATUS_EARLY:INTEGER);
PORT(A:IN STD_LOGIC_VECTOR(C_WIDTH-1 DOWNTO 0);B:IN STD_LOGIC_VECTOR(C_WIDTH-1 DOWNTO 0):=(OTHERS=>'0');OPERATION:IN
 STD_LOGIC_VECTOR(FLT_PT_OPERATION_WIDTH-1 DOWNTO 0);OPERATION_ND:IN STD_LOGIC;OPERATION_RFD:OUT STD_LOGIC;CLK:IN STD_LOGIC;SCLR:IN
 STD_LOGIC;RESULT:OUT STD_LOGIC_VECTOR(C_WIDTH-1 DOWNTO 0);STATUS:OUT STD_LOGIC_VECTOR(FLT_PT_STATUS_WIDTH-1 DOWNTO 0);EXCEPTION:OUT
 STD_LOGIC;UNDERFLOW:OUT STD_LOGIC;OVERFLOW:OUT STD_LOGIC;INVALID_OP:OUT STD_LOGIC;INEXACT:OUT STD_LOGIC;DIVIDE_BY_ZERO:OUT
 STD_LOGIC;DENORM:OUT STD_LOGIC;RDY:OUT STD_LOGIC);END COMPONENT;FUNCTION IIl111Il0IIlOIO000I01l00l0111IIIII(II1111O0III10O0OOlOlOO1l1I1l0IIIII,III00011101l1O1OOI0l0Il0l1l10IIIII:
INTEGER)RETURN INTEGER IS BEGIN IF(II1111O0III10O0OOlOlOO1l1I1l0IIIII=FLT_PT_YES)OR(III00011101l1O1OOI0l0Il0l1l10IIIII=FLT_PT_YES)THEN RETURN(FLT_PT_YES);ELSE RETURN(FLT_PT_NO);
END IF;END;FUNCTION IO0lll11llOIOOIOI1lOOIOl000I0IIIII(IO00OO00lIlIO00llOIll10l0ll1OIIIII:STD_LOGIC_VECTOR(FLT_PT_OPERATION_WIDTH-1 DOWNTO 0))RETURN STD_LOGIC IS BEGIN
 RETURN(IO00OO00lIlIO00llOIll10l0ll1OIIIII(0));END;FUNCTION IIO1lO000Il1O0lOII1IO0OOOIO00IIIII(II1001l0I11O0IIOIl01I1ll0O0OlIIIII:STRING;II1II1OO1ll10IlO0I10O0OI000IIOIIII,IOOl01OO110II1I0lIlI001II11I0IIIII:INTEGER)RETURN STRING IS BEGIN IF(
II1II1OO1ll10IlO0I10O0OI000IIOIIII=FLT_PT_YES)AND(IOOl01OO110II1I0lIlI001II11I0IIIII>=FLT_PT_IS_VIRTEX4)THEN RETURN("virtex4");ELSE RETURN(II1001l0I11O0IIOIl01I1ll0O0OlIIIII);END IF;END;FUNCTION
 II0IIlIOII0IIl1lIO1llO1O1lOlIIIIII(IIll0I0ll1ll1O0IOlO1O01llII00IIIII:STRING;II1ll1Il1Il11O10OllIl0l1l1l0IOIIII,III0II00l1IIlIO100l00OlI1l1O0IIIII:INTEGER)RETURN INTEGER IS BEGIN IF(II1ll1Il1Il11O10OllIl0l1l1l0IOIIII=FLT_PT_YES)AND(
III0II00l1IIlIO100l00OlI1l1O0IIIII>=FLT_PT_IS_VIRTEX4)THEN RETURN(III0II00l1IIlIO100l00OlI1l1O0IIIII-FLT_PT_IS_VIRTEX4);ELSE RETURN(III0II00l1IIlIO100l00OlI1l1O0IIIII);END IF;END;CONSTANT II11OIIIO0I0OI0IIIIO1lOO011IlIIIII:BOOLEAN:=
FLOATING_POINT_V1_0_CHECK(C_FAMILY=>C_FAMILY,C_HAS_ADD=>C_HAS_ADD,C_HAS_SUBTRACT=>C_HAS_SUBTRACT,C_HAS_MULTIPLY=>C_HAS_MULTIPLY,
C_HAS_DIVIDE=>C_HAS_DIVIDE,C_HAS_SQRT=>C_HAS_SQRT,C_HAS_COMPARE=>C_HAS_COMPARE,C_RESULT_WIDTH=>C_RESULT_WIDTH,
C_RESULT_FRACTION_WIDTH=>C_RESULT_FRACTION_WIDTH,C_COMPARE_OPERATION=>C_COMPARE_OPERATION,C_OPTIMIZATION=>C_OPTIMIZATION,
C_MULT_USAGE=>C_MULT_USAGE,C_HAS_SCLR=>C_HAS_SCLR,C_HAS_OPERATION_ND=>C_HAS_OPERATION_ND,C_HAS_OPERATION_RFD=>C_HAS_OPERATION_RFD,
C_HAS_RDY=>C_HAS_RDY,C_HAS_UNDERFLOW=>C_HAS_UNDERFLOW,C_HAS_OVERFLOW=>C_HAS_OVERFLOW,C_HAS_INVALID_OP=>C_HAS_INVALID_OP,
C_HAS_DIVIDE_BY_ZERO=>C_HAS_DIVIDE_BY_ZERO,C_HAS_EXCEPTION=>C_HAS_EXCEPTION,C_STATUS_EARLY=>C_STATUS_EARLY);CONSTANT
 IOl0lI0l0O1IlOIlI1IlO1l01Il00IIIII:INTEGER:=IIl111Il0IIlOIO000I01l00l0111IIIII(C_HAS_ADD,C_HAS_SUBTRACT);CONSTANT III101l00lllOOOlIO0OO1lI1OO1OIIIII:INTEGER:=
FLT_PT_NUMBER_OF_OPERATIONS(C_HAS_ADD,C_HAS_SUBTRACT,C_HAS_MULTIPLY,C_HAS_DIVIDE,C_HAS_SQRT,C_HAS_COMPARE,FLT_PT_NO,FLT_PT_NO);
CONSTANT II0l0l0II0Il010II1l000011O1lIIIIII:BOOLEAN:=(C_HAS_ADD=FLT_PT_YES AND C_HAS_SUBTRACT=FLT_PT_YES);CONSTANT IIlIIOOI1lOO0O0I1O1O10lI0OlIOOIIII:STRING:=
IIO1lO000Il1O0lOII1IO0OOOIO00IIIII(C_FAMILY,C_HAS_MULTIPLY,C_MULT_USAGE);CONSTANT IOO0lOOOll1OI0OI0lI10IOOOII00IIIII:INTEGER:=II0IIlIOII0IIl1lIO1llO1O1lOlIIIIII(C_FAMILY,
C_HAS_MULTIPLY,C_MULT_USAGE);SIGNAL II111O1llOOlI0lOOIIIl0OIlIlllIIIII:STD_LOGIC;SIGNAL IIO11lIl110IO0lO00IOOl0Il11I1IIIII:STD_LOGIC;SIGNAL II1IO0OO0IOlO11110OOlO1O0101IOIIII:STD_LOGIC;SIGNAL
 II0lIlIIOl0I0Ol0lIl0111l1I1l1IIIII:STD_LOGIC;SIGNAL IO0OIl1OO10lO00IlIl0Il0l1l1OIIIIII:STD_LOGIC;SIGNAL IO0lllOII000O01100OOI0II1II01IIIII:STD_LOGIC;SIGNAL IO0IllIIO11IlI1010IIl0l000001IIIII:STD_LOGIC;SIGNAL II1l0I0l10l0I1I1lO01l10I01lI1IIIII:
STD_LOGIC;SIGNAL IIO001lIl0II1lI10I1000O00Ol10IIIII:STD_LOGIC_VECTOR(FLT_PT_STATUS_WIDTH-1 DOWNTO 0);SIGNAL IIOI1lO0I00III00II0IO0ll0111IOIIII:STD_LOGIC;SIGNAL III11OII1IlIl1001I1IO1111l0IlIIIII:
STD_LOGIC_VECTOR(FLT_PT_OPERATION_WIDTH-1 DOWNTO 0);BEGIN YES_SCLR:IF C_HAS_SCLR=FLT_PT_YES GENERATE IO0OIl1OO10lO00IlIl0Il0l1l1OIIIIII<=SCLR;END GENERATE;
NO_SCLR:IF C_HAS_SCLR/=FLT_PT_YES GENERATE IO0OIl1OO10lO00IlIl0Il0l1l1OIIIIII<='0';END GENERATE;YES_OPERATION_ND:IF C_HAS_OPERATION_ND=FLT_PT_YES GENERATE
 IO0lllOII000O01100OOI0II1II01IIIII<=OPERATION_ND;END GENERATE;NO_OPERATION_ND:IF C_HAS_OPERATION_ND/=FLT_PT_YES GENERATE IO0lllOII000O01100OOI0II1II01IIIII<='1';END
 GENERATE;YES_OPERATION_RFD:IF C_HAS_OPERATION_RFD=FLT_PT_YES GENERATE OPERATION_RFD<=IO0IllIIO11IlI1010IIl0l000001IIIII;END GENERATE;NO_OPERATION_RFD
:IF C_HAS_OPERATION_RFD/=FLT_PT_YES GENERATE OPERATION_RFD<='X';END GENERATE;YES_RDY:IF C_HAS_RDY=FLT_PT_YES GENERATE RDY<=II1l0I0l10l0I1I1lO01l10I01lI1IIIII;
END GENERATE;NO_RDY:IF C_HAS_RDY/=FLT_PT_YES GENERATE RDY<='X';END GENERATE;YES_UNDERFLOW:IF C_HAS_UNDERFLOW=FLT_PT_YES GENERATE
 UNDERFLOW<=II111O1llOOlI0lOOIIIl0OIlIlllIIIII;END GENERATE;NO_UNDERFLOW:IF C_HAS_UNDERFLOW/=FLT_PT_YES GENERATE UNDERFLOW<='X';END GENERATE;YES_OVERFLOW
:IF C_HAS_OVERFLOW=FLT_PT_YES GENERATE OVERFLOW<=IIO11lIl110IO0lO00IOOl0Il11I1IIIII;END GENERATE;NO_OVERFLOW:IF C_HAS_OVERFLOW/=FLT_PT_YES GENERATE
 OVERFLOW<='X';END GENERATE;YES_INVALID_OP:IF C_HAS_INVALID_OP=FLT_PT_YES GENERATE INVALID_OP<=II0lIlIIOl0I0Ol0lIl0111l1I1l1IIIII;END GENERATE;
NO_INVALID_OP:IF C_HAS_INVALID_OP/=FLT_PT_YES GENERATE INVALID_OP<='X';END GENERATE;YES_DIVIDE_BY_ZERO:IF(C_HAS_DIVIDE_BY_ZERO=
FLT_PT_YES)GENERATE DIVIDE_BY_ZERO<=II1IO0OO0IOlO11110OOlO1O0101IOIIII;END GENERATE;NO_DIVIDE_BY_ZERO:IF(C_HAS_DIVIDE_BY_ZERO/=FLT_PT_YES)GENERATE
 DIVIDE_BY_ZERO<='X';END GENERATE;YES_EXCEPTION:IF C_HAS_EXCEPTION=FLT_PT_YES GENERATE EXCEPTION<=IIOI1lO0I00III00II0IO0ll0111IOIIII;END GENERATE;
NO_EXCEPTION:IF C_HAS_EXCEPTION/=FLT_PT_YES GENERATE EXCEPTION<='X';END GENERATE;YES_STATUS:IF C_HAS_STATUS=FLT_PT_YES GENERATE
 STATUS<=IIO001lIl0II1lI10I1000O00Ol10IIIII;END GENERATE;NO_STATUS:IF C_HAS_STATUS=FLT_PT_NO GENERATE STATUS<=(OTHERS=>'X');END GENERATE;YES_COMPARE:IF
 C_HAS_COMPARE=FLT_PT_YES GENERATE PROG_COMPARE:IF C_COMPARE_OPERATION=FLT_PT_PROGRAMMABLE GENERATE III11OII1IlIl1001I1IO1111l0IlIIIII(
FLT_PT_COMPARE_OPERATION_SLICE)<=OPERATION(FLT_PT_COMPARE_OPERATION_SLICE);END GENERATE;FIXED_COMPARE:IF C_COMPARE_OPERATION/=
FLT_PT_PROGRAMMABLE GENERATE III11OII1IlIl1001I1IO1111l0IlIIIII(FLT_PT_COMPARE_OPERATION_SLICE)<=STD_LOGIC_VECTOR(TO_UNSIGNED(C_COMPARE_OPERATION,
FLT_PT_COMPARE_OPERATION_WIDTH));END GENERATE;END GENERATE;OPERATION_RQD:IF III101l00lllOOOlIO0OO1lI1OO1OIIIII>1 GENERATE III11OII1IlIl1001I1IO1111l0IlIIIII(
FLT_PT_OP_CODE_SLICE)<=OPERATION(FLT_PT_OP_CODE_SLICE);END GENERATE;ONE_OPERATION:IF III101l00lllOOOlIO0OO1lI1OO1OIIIII=1 GENERATE CONSTANT
 IIII11lI1lOl0OlOO0II11lI101lOIIIII:STD_LOGIC_VECTOR(FLT_PT_OP_CODE_SLICE):=FLT_PT_GET_OP_CODE(C_HAS_ADD,C_HAS_SUBTRACT,C_HAS_MULTIPLY,C_HAS_DIVIDE,
C_HAS_SQRT,C_HAS_COMPARE,C_HAS_FIX_TO_FLT,C_HAS_FLT_TO_FIX);BEGIN III11OII1IlIl1001I1IO1111l0IlIIIII(FLT_PT_OP_CODE_SLICE)<=IIII11lI1lOl0OlOO0II11lI101lOIIIII;END GENERATE;
FP_OP:FLT_PT_OPERATOR GENERIC MAP(C_FAMILY=>IIlIIOOI1lOO0O0I1O1O10lI0OlIOOIIII,C_WIDTH=>C_RESULT_WIDTH,C_FRACTION_WIDTH=>C_RESULT_FRACTION_WIDTH,
C_OPTIMIZATION=>C_OPTIMIZATION,C_MULT_USAGE=>IOO0lOOOll1OI0OI0lI10IOOOII00IIIII,C_HAS_STATUS=>C_HAS_STATUS,C_STATUS_EARLY=>C_STATUS_EARLY)PORT MAP(A
=>A,B=>B,OPERATION=>III11OII1IlIl1001I1IO1111l0IlIIIII,OPERATION_ND=>IO0lllOII000O01100OOI0II1II01IIIII,OPERATION_RFD=>IO0IllIIO11IlI1010IIl0l000001IIIII,CLK=>CLK,SCLR=>IO0OIl1OO10lO00IlIl0Il0l1l1OIIIIII,RESULT=>RESULT
,STATUS=>IIO001lIl0II1lI10I1000O00Ol10IIIII,EXCEPTION=>IIOI1lO0I00III00II0IO0ll0111IOIIII,UNDERFLOW=>II111O1llOOlI0lOOIIIl0OIlIlllIIIII,OVERFLOW=>IIO11lIl110IO0lO00IOOl0Il11I1IIIII,INVALID_OP=>II0lIlIIOl0I0Ol0lIl0111l1I1l1IIIII,DIVIDE_BY_ZERO=>
II1IO0OO0IOlO11110OOlO1O0101IOIIII,RDY=>II1l0I0l10l0I1I1lO01l10I01lI1IIIII);END;
